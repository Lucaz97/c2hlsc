
//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_inout_prereg_en_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2019 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_inout_prereg_en_v1 (din, ldout, dout, zin, lzout, zout);

    parameter integer rscid = 1;
    parameter integer width = 8;

    output [width-1:0] din;
    input              ldout;
    input  [width-1:0] dout;
    input  [width-1:0] zin;
    output             lzout;
    output [width-1:0] zout;

    wire   [width-1:0] din;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzout = ldout;
    assign din = zin;
    assign zout = dout;

endmodule



//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   lc4976@hansolo.poly.edu
//  Generated date: Tue Apr  9 23:24:51 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    MixColumns_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module MixColumns_core_core_fsm (
  clk, rst_n, fsm_output, for_C_1_tr0
);
  input clk;
  input rst_n;
  output [3:0] fsm_output;
  reg [3:0] fsm_output;
  input for_C_1_tr0;


  // FSM State Type Declaration for MixColumns_core_core_fsm_1
  parameter
    main_C_0 = 2'd0,
    for_C_0 = 2'd1,
    for_C_1 = 2'd2,
    main_C_1 = 2'd3;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : MixColumns_core_core_fsm_1
    case (state_var)
      for_C_0 : begin
        fsm_output = 4'b0010;
        state_var_NS = for_C_1;
      end
      for_C_1 : begin
        fsm_output = 4'b0100;
        if ( for_C_1_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 4'b1000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 4'b0001;
        state_var_NS = for_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MixColumns_core
// ------------------------------------------------------------------


module MixColumns_core (
  clk, rst_n, state_rsc_zout, state_rsc_lzout, state_rsc_zin, state_triosy_lz
);
  input clk;
  input rst_n;
  output [127:0] state_rsc_zout;
  output state_rsc_lzout;
  input [127:0] state_rsc_zin;
  output state_triosy_lz;


  // Interconnect Declarations
  wire [127:0] state_rsci_din;
  reg state_triosy_obj_ld;
  wire [3:0] fsm_output;
  wire and_dcpl;
  wire or_dcpl_1;
  wire or_dcpl_2;
  wire or_dcpl_3;
  wire [2:0] i_2_0_sva_2;
  wire [3:0] nl_i_2_0_sva_2;
  reg [1:0] i_2_0_sva_1_0;
  wire for_conc_35_cmx_7_sva_1;
  wire for_conc_35_cmx_6_sva_1;
  wire for_conc_35_cmx_5_sva_1;
  wire for_conc_35_cmx_4_sva_1;
  wire for_conc_35_cmx_3_sva_1;
  wire for_conc_35_cmx_2_sva_1;
  wire for_conc_35_cmx_1_sva_1;
  wire for_conc_35_cmx_0_sva_1;
  wire for_conc_34_cmx_7_sva_1;
  wire for_conc_34_cmx_6_sva_1;
  wire for_conc_34_cmx_5_sva_1;
  wire for_conc_34_cmx_4_sva_1;
  wire for_conc_34_cmx_3_sva_1;
  wire for_conc_34_cmx_2_sva_1;
  wire for_conc_34_cmx_1_sva_1;
  wire for_conc_34_cmx_0_sva_1;
  wire for_conc_33_cmx_7_sva_1;
  wire for_conc_33_cmx_6_sva_1;
  wire for_conc_33_cmx_5_sva_1;
  wire for_conc_33_cmx_4_sva_1;
  wire for_conc_33_cmx_3_sva_1;
  wire for_conc_33_cmx_2_sva_1;
  wire for_conc_33_cmx_1_sva_1;
  wire for_conc_33_cmx_0_sva_1;
  wire for_conc_32_cmx_7_sva_1;
  wire for_conc_32_cmx_6_sva_1;
  wire for_conc_32_cmx_5_sva_1;
  wire for_conc_32_cmx_4_sva_1;
  wire for_conc_32_cmx_3_sva_1;
  wire for_conc_32_cmx_2_sva_1;
  wire for_conc_32_cmx_1_sva_1;
  wire for_conc_32_cmx_0_sva_1;
  wire [7:0] for_slc_state_8_7_0_4_ncse_sva_1;
  wire [7:0] t_sva_1;
  wire [7:0] Tmp_sva_1;
  wire [7:0] for_slc_state_8_7_0_3_ncse_sva_1;
  wire [7:0] for_slc_state_8_7_0_2_cse_sva_1;
  wire xor_cse;
  wire xor_cse_1;
  wire xor_cse_2;
  wire xor_cse_3;
  wire xor_cse_4;
  wire xor_cse_5;

  wire i_not_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_state_rsci_ldout;
  assign nl_state_rsci_ldout = fsm_output[1];
  wire for_mux_127_nl;
  wire for_mux_126_nl;
  wire for_mux_125_nl;
  wire for_mux_124_nl;
  wire for_mux_123_nl;
  wire for_mux_122_nl;
  wire for_mux_121_nl;
  wire for_mux_120_nl;
  wire for_mux_119_nl;
  wire for_mux_118_nl;
  wire for_mux_117_nl;
  wire for_mux_116_nl;
  wire for_mux_115_nl;
  wire for_mux_114_nl;
  wire for_mux_113_nl;
  wire for_mux_112_nl;
  wire for_mux_111_nl;
  wire for_mux_110_nl;
  wire for_mux_109_nl;
  wire for_mux_108_nl;
  wire for_mux_107_nl;
  wire for_mux_106_nl;
  wire for_mux_105_nl;
  wire for_mux_104_nl;
  wire for_mux_103_nl;
  wire for_mux_102_nl;
  wire for_mux_101_nl;
  wire for_mux_100_nl;
  wire for_mux_99_nl;
  wire for_mux_98_nl;
  wire for_mux_97_nl;
  wire for_mux_96_nl;
  wire for_mux_95_nl;
  wire for_mux_94_nl;
  wire for_mux_93_nl;
  wire for_mux_92_nl;
  wire for_mux_91_nl;
  wire for_mux_90_nl;
  wire for_mux_89_nl;
  wire for_mux_88_nl;
  wire for_mux_87_nl;
  wire for_mux_86_nl;
  wire for_mux_85_nl;
  wire for_mux_84_nl;
  wire for_mux_83_nl;
  wire for_mux_82_nl;
  wire for_mux_81_nl;
  wire for_mux_80_nl;
  wire for_mux_79_nl;
  wire for_mux_78_nl;
  wire for_mux_77_nl;
  wire for_mux_76_nl;
  wire for_mux_75_nl;
  wire for_mux_74_nl;
  wire for_mux_73_nl;
  wire for_mux_72_nl;
  wire for_mux_71_nl;
  wire for_mux_70_nl;
  wire for_mux_69_nl;
  wire for_mux_68_nl;
  wire for_mux_67_nl;
  wire for_mux_66_nl;
  wire for_mux_65_nl;
  wire for_mux_64_nl;
  wire for_mux_63_nl;
  wire for_mux_62_nl;
  wire for_mux_61_nl;
  wire for_mux_60_nl;
  wire for_mux_59_nl;
  wire for_mux_58_nl;
  wire for_mux_57_nl;
  wire for_mux_56_nl;
  wire for_mux_55_nl;
  wire for_mux_54_nl;
  wire for_mux_53_nl;
  wire for_mux_52_nl;
  wire for_mux_51_nl;
  wire for_mux_50_nl;
  wire for_mux_49_nl;
  wire for_mux_48_nl;
  wire for_mux_47_nl;
  wire for_mux_46_nl;
  wire for_mux_45_nl;
  wire for_mux_44_nl;
  wire for_mux_43_nl;
  wire for_mux_42_nl;
  wire for_mux_41_nl;
  wire for_mux_40_nl;
  wire for_mux_39_nl;
  wire for_mux_38_nl;
  wire for_mux_37_nl;
  wire for_mux_36_nl;
  wire for_mux_35_nl;
  wire for_mux_34_nl;
  wire for_mux_33_nl;
  wire for_mux_32_nl;
  wire for_mux_31_nl;
  wire for_mux_30_nl;
  wire for_mux_29_nl;
  wire for_mux_28_nl;
  wire for_mux_27_nl;
  wire for_mux_26_nl;
  wire for_mux_25_nl;
  wire for_mux_24_nl;
  wire for_mux_23_nl;
  wire for_mux_22_nl;
  wire for_mux_21_nl;
  wire for_mux_20_nl;
  wire for_mux_19_nl;
  wire for_mux_18_nl;
  wire for_mux_17_nl;
  wire for_mux_16_nl;
  wire for_mux_15_nl;
  wire for_mux_14_nl;
  wire for_mux_13_nl;
  wire for_mux_12_nl;
  wire for_mux_11_nl;
  wire for_mux_10_nl;
  wire for_mux_9_nl;
  wire for_mux_8_nl;
  wire for_mux_7_nl;
  wire for_mux_6_nl;
  wire for_mux_5_nl;
  wire for_mux_4_nl;
  wire for_mux_3_nl;
  wire for_mux_2_nl;
  wire for_mux_1_nl;
  wire for_mux_nl;
  wire [127:0] nl_state_rsci_dout;
  assign for_mux_127_nl = MUX_s_1_2_2(for_conc_35_cmx_7_sva_1, (state_rsci_din[127]),
      or_dcpl_3);
  assign for_mux_126_nl = MUX_s_1_2_2(for_conc_35_cmx_6_sva_1, (state_rsci_din[126]),
      or_dcpl_3);
  assign for_mux_125_nl = MUX_s_1_2_2(for_conc_35_cmx_5_sva_1, (state_rsci_din[125]),
      or_dcpl_3);
  assign for_mux_124_nl = MUX_s_1_2_2(for_conc_35_cmx_4_sva_1, (state_rsci_din[124]),
      or_dcpl_3);
  assign for_mux_123_nl = MUX_s_1_2_2(for_conc_35_cmx_3_sva_1, (state_rsci_din[123]),
      or_dcpl_3);
  assign for_mux_122_nl = MUX_s_1_2_2(for_conc_35_cmx_2_sva_1, (state_rsci_din[122]),
      or_dcpl_3);
  assign for_mux_121_nl = MUX_s_1_2_2(for_conc_35_cmx_1_sva_1, (state_rsci_din[121]),
      or_dcpl_3);
  assign for_mux_120_nl = MUX_s_1_2_2(for_conc_35_cmx_0_sva_1, (state_rsci_din[120]),
      or_dcpl_3);
  assign for_mux_119_nl = MUX_s_1_2_2(for_conc_34_cmx_7_sva_1, (state_rsci_din[119]),
      or_dcpl_3);
  assign for_mux_118_nl = MUX_s_1_2_2(for_conc_34_cmx_6_sva_1, (state_rsci_din[118]),
      or_dcpl_3);
  assign for_mux_117_nl = MUX_s_1_2_2(for_conc_34_cmx_5_sva_1, (state_rsci_din[117]),
      or_dcpl_3);
  assign for_mux_116_nl = MUX_s_1_2_2(for_conc_34_cmx_4_sva_1, (state_rsci_din[116]),
      or_dcpl_3);
  assign for_mux_115_nl = MUX_s_1_2_2(for_conc_34_cmx_3_sva_1, (state_rsci_din[115]),
      or_dcpl_3);
  assign for_mux_114_nl = MUX_s_1_2_2(for_conc_34_cmx_2_sva_1, (state_rsci_din[114]),
      or_dcpl_3);
  assign for_mux_113_nl = MUX_s_1_2_2(for_conc_34_cmx_1_sva_1, (state_rsci_din[113]),
      or_dcpl_3);
  assign for_mux_112_nl = MUX_s_1_2_2(for_conc_34_cmx_0_sva_1, (state_rsci_din[112]),
      or_dcpl_3);
  assign for_mux_111_nl = MUX_s_1_2_2(for_conc_33_cmx_7_sva_1, (state_rsci_din[111]),
      or_dcpl_3);
  assign for_mux_110_nl = MUX_s_1_2_2(for_conc_33_cmx_6_sva_1, (state_rsci_din[110]),
      or_dcpl_3);
  assign for_mux_109_nl = MUX_s_1_2_2(for_conc_33_cmx_5_sva_1, (state_rsci_din[109]),
      or_dcpl_3);
  assign for_mux_108_nl = MUX_s_1_2_2(for_conc_33_cmx_4_sva_1, (state_rsci_din[108]),
      or_dcpl_3);
  assign for_mux_107_nl = MUX_s_1_2_2(for_conc_33_cmx_3_sva_1, (state_rsci_din[107]),
      or_dcpl_3);
  assign for_mux_106_nl = MUX_s_1_2_2(for_conc_33_cmx_2_sva_1, (state_rsci_din[106]),
      or_dcpl_3);
  assign for_mux_105_nl = MUX_s_1_2_2(for_conc_33_cmx_1_sva_1, (state_rsci_din[105]),
      or_dcpl_3);
  assign for_mux_104_nl = MUX_s_1_2_2(for_conc_33_cmx_0_sva_1, (state_rsci_din[104]),
      or_dcpl_3);
  assign for_mux_103_nl = MUX_s_1_2_2(for_conc_32_cmx_7_sva_1, (state_rsci_din[103]),
      or_dcpl_3);
  assign for_mux_102_nl = MUX_s_1_2_2(for_conc_32_cmx_6_sva_1, (state_rsci_din[102]),
      or_dcpl_3);
  assign for_mux_101_nl = MUX_s_1_2_2(for_conc_32_cmx_5_sva_1, (state_rsci_din[101]),
      or_dcpl_3);
  assign for_mux_100_nl = MUX_s_1_2_2(for_conc_32_cmx_4_sva_1, (state_rsci_din[100]),
      or_dcpl_3);
  assign for_mux_99_nl = MUX_s_1_2_2(for_conc_32_cmx_3_sva_1, (state_rsci_din[99]),
      or_dcpl_3);
  assign for_mux_98_nl = MUX_s_1_2_2(for_conc_32_cmx_2_sva_1, (state_rsci_din[98]),
      or_dcpl_3);
  assign for_mux_97_nl = MUX_s_1_2_2(for_conc_32_cmx_1_sva_1, (state_rsci_din[97]),
      or_dcpl_3);
  assign for_mux_96_nl = MUX_s_1_2_2(for_conc_32_cmx_0_sva_1, (state_rsci_din[96]),
      or_dcpl_3);
  assign for_mux_95_nl = MUX_s_1_2_2(for_conc_35_cmx_7_sva_1, (state_rsci_din[95]),
      or_dcpl_2);
  assign for_mux_94_nl = MUX_s_1_2_2(for_conc_35_cmx_6_sva_1, (state_rsci_din[94]),
      or_dcpl_2);
  assign for_mux_93_nl = MUX_s_1_2_2(for_conc_35_cmx_5_sva_1, (state_rsci_din[93]),
      or_dcpl_2);
  assign for_mux_92_nl = MUX_s_1_2_2(for_conc_35_cmx_4_sva_1, (state_rsci_din[92]),
      or_dcpl_2);
  assign for_mux_91_nl = MUX_s_1_2_2(for_conc_35_cmx_3_sva_1, (state_rsci_din[91]),
      or_dcpl_2);
  assign for_mux_90_nl = MUX_s_1_2_2(for_conc_35_cmx_2_sva_1, (state_rsci_din[90]),
      or_dcpl_2);
  assign for_mux_89_nl = MUX_s_1_2_2(for_conc_35_cmx_1_sva_1, (state_rsci_din[89]),
      or_dcpl_2);
  assign for_mux_88_nl = MUX_s_1_2_2(for_conc_35_cmx_0_sva_1, (state_rsci_din[88]),
      or_dcpl_2);
  assign for_mux_87_nl = MUX_s_1_2_2(for_conc_34_cmx_7_sva_1, (state_rsci_din[87]),
      or_dcpl_2);
  assign for_mux_86_nl = MUX_s_1_2_2(for_conc_34_cmx_6_sva_1, (state_rsci_din[86]),
      or_dcpl_2);
  assign for_mux_85_nl = MUX_s_1_2_2(for_conc_34_cmx_5_sva_1, (state_rsci_din[85]),
      or_dcpl_2);
  assign for_mux_84_nl = MUX_s_1_2_2(for_conc_34_cmx_4_sva_1, (state_rsci_din[84]),
      or_dcpl_2);
  assign for_mux_83_nl = MUX_s_1_2_2(for_conc_34_cmx_3_sva_1, (state_rsci_din[83]),
      or_dcpl_2);
  assign for_mux_82_nl = MUX_s_1_2_2(for_conc_34_cmx_2_sva_1, (state_rsci_din[82]),
      or_dcpl_2);
  assign for_mux_81_nl = MUX_s_1_2_2(for_conc_34_cmx_1_sva_1, (state_rsci_din[81]),
      or_dcpl_2);
  assign for_mux_80_nl = MUX_s_1_2_2(for_conc_34_cmx_0_sva_1, (state_rsci_din[80]),
      or_dcpl_2);
  assign for_mux_79_nl = MUX_s_1_2_2(for_conc_33_cmx_7_sva_1, (state_rsci_din[79]),
      or_dcpl_2);
  assign for_mux_78_nl = MUX_s_1_2_2(for_conc_33_cmx_6_sva_1, (state_rsci_din[78]),
      or_dcpl_2);
  assign for_mux_77_nl = MUX_s_1_2_2(for_conc_33_cmx_5_sva_1, (state_rsci_din[77]),
      or_dcpl_2);
  assign for_mux_76_nl = MUX_s_1_2_2(for_conc_33_cmx_4_sva_1, (state_rsci_din[76]),
      or_dcpl_2);
  assign for_mux_75_nl = MUX_s_1_2_2(for_conc_33_cmx_3_sva_1, (state_rsci_din[75]),
      or_dcpl_2);
  assign for_mux_74_nl = MUX_s_1_2_2(for_conc_33_cmx_2_sva_1, (state_rsci_din[74]),
      or_dcpl_2);
  assign for_mux_73_nl = MUX_s_1_2_2(for_conc_33_cmx_1_sva_1, (state_rsci_din[73]),
      or_dcpl_2);
  assign for_mux_72_nl = MUX_s_1_2_2(for_conc_33_cmx_0_sva_1, (state_rsci_din[72]),
      or_dcpl_2);
  assign for_mux_71_nl = MUX_s_1_2_2(for_conc_32_cmx_7_sva_1, (state_rsci_din[71]),
      or_dcpl_2);
  assign for_mux_70_nl = MUX_s_1_2_2(for_conc_32_cmx_6_sva_1, (state_rsci_din[70]),
      or_dcpl_2);
  assign for_mux_69_nl = MUX_s_1_2_2(for_conc_32_cmx_5_sva_1, (state_rsci_din[69]),
      or_dcpl_2);
  assign for_mux_68_nl = MUX_s_1_2_2(for_conc_32_cmx_4_sva_1, (state_rsci_din[68]),
      or_dcpl_2);
  assign for_mux_67_nl = MUX_s_1_2_2(for_conc_32_cmx_3_sva_1, (state_rsci_din[67]),
      or_dcpl_2);
  assign for_mux_66_nl = MUX_s_1_2_2(for_conc_32_cmx_2_sva_1, (state_rsci_din[66]),
      or_dcpl_2);
  assign for_mux_65_nl = MUX_s_1_2_2(for_conc_32_cmx_1_sva_1, (state_rsci_din[65]),
      or_dcpl_2);
  assign for_mux_64_nl = MUX_s_1_2_2(for_conc_32_cmx_0_sva_1, (state_rsci_din[64]),
      or_dcpl_2);
  assign for_mux_63_nl = MUX_s_1_2_2(for_conc_35_cmx_7_sva_1, (state_rsci_din[63]),
      or_dcpl_1);
  assign for_mux_62_nl = MUX_s_1_2_2(for_conc_35_cmx_6_sva_1, (state_rsci_din[62]),
      or_dcpl_1);
  assign for_mux_61_nl = MUX_s_1_2_2(for_conc_35_cmx_5_sva_1, (state_rsci_din[61]),
      or_dcpl_1);
  assign for_mux_60_nl = MUX_s_1_2_2(for_conc_35_cmx_4_sva_1, (state_rsci_din[60]),
      or_dcpl_1);
  assign for_mux_59_nl = MUX_s_1_2_2(for_conc_35_cmx_3_sva_1, (state_rsci_din[59]),
      or_dcpl_1);
  assign for_mux_58_nl = MUX_s_1_2_2(for_conc_35_cmx_2_sva_1, (state_rsci_din[58]),
      or_dcpl_1);
  assign for_mux_57_nl = MUX_s_1_2_2(for_conc_35_cmx_1_sva_1, (state_rsci_din[57]),
      or_dcpl_1);
  assign for_mux_56_nl = MUX_s_1_2_2(for_conc_35_cmx_0_sva_1, (state_rsci_din[56]),
      or_dcpl_1);
  assign for_mux_55_nl = MUX_s_1_2_2(for_conc_34_cmx_7_sva_1, (state_rsci_din[55]),
      or_dcpl_1);
  assign for_mux_54_nl = MUX_s_1_2_2(for_conc_34_cmx_6_sva_1, (state_rsci_din[54]),
      or_dcpl_1);
  assign for_mux_53_nl = MUX_s_1_2_2(for_conc_34_cmx_5_sva_1, (state_rsci_din[53]),
      or_dcpl_1);
  assign for_mux_52_nl = MUX_s_1_2_2(for_conc_34_cmx_4_sva_1, (state_rsci_din[52]),
      or_dcpl_1);
  assign for_mux_51_nl = MUX_s_1_2_2(for_conc_34_cmx_3_sva_1, (state_rsci_din[51]),
      or_dcpl_1);
  assign for_mux_50_nl = MUX_s_1_2_2(for_conc_34_cmx_2_sva_1, (state_rsci_din[50]),
      or_dcpl_1);
  assign for_mux_49_nl = MUX_s_1_2_2(for_conc_34_cmx_1_sva_1, (state_rsci_din[49]),
      or_dcpl_1);
  assign for_mux_48_nl = MUX_s_1_2_2(for_conc_34_cmx_0_sva_1, (state_rsci_din[48]),
      or_dcpl_1);
  assign for_mux_47_nl = MUX_s_1_2_2(for_conc_33_cmx_7_sva_1, (state_rsci_din[47]),
      or_dcpl_1);
  assign for_mux_46_nl = MUX_s_1_2_2(for_conc_33_cmx_6_sva_1, (state_rsci_din[46]),
      or_dcpl_1);
  assign for_mux_45_nl = MUX_s_1_2_2(for_conc_33_cmx_5_sva_1, (state_rsci_din[45]),
      or_dcpl_1);
  assign for_mux_44_nl = MUX_s_1_2_2(for_conc_33_cmx_4_sva_1, (state_rsci_din[44]),
      or_dcpl_1);
  assign for_mux_43_nl = MUX_s_1_2_2(for_conc_33_cmx_3_sva_1, (state_rsci_din[43]),
      or_dcpl_1);
  assign for_mux_42_nl = MUX_s_1_2_2(for_conc_33_cmx_2_sva_1, (state_rsci_din[42]),
      or_dcpl_1);
  assign for_mux_41_nl = MUX_s_1_2_2(for_conc_33_cmx_1_sva_1, (state_rsci_din[41]),
      or_dcpl_1);
  assign for_mux_40_nl = MUX_s_1_2_2(for_conc_33_cmx_0_sva_1, (state_rsci_din[40]),
      or_dcpl_1);
  assign for_mux_39_nl = MUX_s_1_2_2(for_conc_32_cmx_7_sva_1, (state_rsci_din[39]),
      or_dcpl_1);
  assign for_mux_38_nl = MUX_s_1_2_2(for_conc_32_cmx_6_sva_1, (state_rsci_din[38]),
      or_dcpl_1);
  assign for_mux_37_nl = MUX_s_1_2_2(for_conc_32_cmx_5_sva_1, (state_rsci_din[37]),
      or_dcpl_1);
  assign for_mux_36_nl = MUX_s_1_2_2(for_conc_32_cmx_4_sva_1, (state_rsci_din[36]),
      or_dcpl_1);
  assign for_mux_35_nl = MUX_s_1_2_2(for_conc_32_cmx_3_sva_1, (state_rsci_din[35]),
      or_dcpl_1);
  assign for_mux_34_nl = MUX_s_1_2_2(for_conc_32_cmx_2_sva_1, (state_rsci_din[34]),
      or_dcpl_1);
  assign for_mux_33_nl = MUX_s_1_2_2(for_conc_32_cmx_1_sva_1, (state_rsci_din[33]),
      or_dcpl_1);
  assign for_mux_32_nl = MUX_s_1_2_2(for_conc_32_cmx_0_sva_1, (state_rsci_din[32]),
      or_dcpl_1);
  assign for_mux_31_nl = MUX_s_1_2_2((state_rsci_din[31]), for_conc_35_cmx_7_sva_1,
      and_dcpl);
  assign for_mux_30_nl = MUX_s_1_2_2((state_rsci_din[30]), for_conc_35_cmx_6_sva_1,
      and_dcpl);
  assign for_mux_29_nl = MUX_s_1_2_2((state_rsci_din[29]), for_conc_35_cmx_5_sva_1,
      and_dcpl);
  assign for_mux_28_nl = MUX_s_1_2_2((state_rsci_din[28]), for_conc_35_cmx_4_sva_1,
      and_dcpl);
  assign for_mux_27_nl = MUX_s_1_2_2((state_rsci_din[27]), for_conc_35_cmx_3_sva_1,
      and_dcpl);
  assign for_mux_26_nl = MUX_s_1_2_2((state_rsci_din[26]), for_conc_35_cmx_2_sva_1,
      and_dcpl);
  assign for_mux_25_nl = MUX_s_1_2_2((state_rsci_din[25]), for_conc_35_cmx_1_sva_1,
      and_dcpl);
  assign for_mux_24_nl = MUX_s_1_2_2((state_rsci_din[24]), for_conc_35_cmx_0_sva_1,
      and_dcpl);
  assign for_mux_23_nl = MUX_s_1_2_2((state_rsci_din[23]), for_conc_34_cmx_7_sva_1,
      and_dcpl);
  assign for_mux_22_nl = MUX_s_1_2_2((state_rsci_din[22]), for_conc_34_cmx_6_sva_1,
      and_dcpl);
  assign for_mux_21_nl = MUX_s_1_2_2((state_rsci_din[21]), for_conc_34_cmx_5_sva_1,
      and_dcpl);
  assign for_mux_20_nl = MUX_s_1_2_2((state_rsci_din[20]), for_conc_34_cmx_4_sva_1,
      and_dcpl);
  assign for_mux_19_nl = MUX_s_1_2_2((state_rsci_din[19]), for_conc_34_cmx_3_sva_1,
      and_dcpl);
  assign for_mux_18_nl = MUX_s_1_2_2((state_rsci_din[18]), for_conc_34_cmx_2_sva_1,
      and_dcpl);
  assign for_mux_17_nl = MUX_s_1_2_2((state_rsci_din[17]), for_conc_34_cmx_1_sva_1,
      and_dcpl);
  assign for_mux_16_nl = MUX_s_1_2_2((state_rsci_din[16]), for_conc_34_cmx_0_sva_1,
      and_dcpl);
  assign for_mux_15_nl = MUX_s_1_2_2((state_rsci_din[15]), for_conc_33_cmx_7_sva_1,
      and_dcpl);
  assign for_mux_14_nl = MUX_s_1_2_2((state_rsci_din[14]), for_conc_33_cmx_6_sva_1,
      and_dcpl);
  assign for_mux_13_nl = MUX_s_1_2_2((state_rsci_din[13]), for_conc_33_cmx_5_sva_1,
      and_dcpl);
  assign for_mux_12_nl = MUX_s_1_2_2((state_rsci_din[12]), for_conc_33_cmx_4_sva_1,
      and_dcpl);
  assign for_mux_11_nl = MUX_s_1_2_2((state_rsci_din[11]), for_conc_33_cmx_3_sva_1,
      and_dcpl);
  assign for_mux_10_nl = MUX_s_1_2_2((state_rsci_din[10]), for_conc_33_cmx_2_sva_1,
      and_dcpl);
  assign for_mux_9_nl = MUX_s_1_2_2((state_rsci_din[9]), for_conc_33_cmx_1_sva_1,
      and_dcpl);
  assign for_mux_8_nl = MUX_s_1_2_2((state_rsci_din[8]), for_conc_33_cmx_0_sva_1,
      and_dcpl);
  assign for_mux_7_nl = MUX_s_1_2_2((state_rsci_din[7]), for_conc_32_cmx_7_sva_1,
      and_dcpl);
  assign for_mux_6_nl = MUX_s_1_2_2((state_rsci_din[6]), for_conc_32_cmx_6_sva_1,
      and_dcpl);
  assign for_mux_5_nl = MUX_s_1_2_2((state_rsci_din[5]), for_conc_32_cmx_5_sva_1,
      and_dcpl);
  assign for_mux_4_nl = MUX_s_1_2_2((state_rsci_din[4]), for_conc_32_cmx_4_sva_1,
      and_dcpl);
  assign for_mux_3_nl = MUX_s_1_2_2((state_rsci_din[3]), for_conc_32_cmx_3_sva_1,
      and_dcpl);
  assign for_mux_2_nl = MUX_s_1_2_2((state_rsci_din[2]), for_conc_32_cmx_2_sva_1,
      and_dcpl);
  assign for_mux_1_nl = MUX_s_1_2_2((state_rsci_din[1]), for_conc_32_cmx_1_sva_1,
      and_dcpl);
  assign for_mux_nl = MUX_s_1_2_2((state_rsci_din[0]), for_conc_32_cmx_0_sva_1, and_dcpl);
  assign nl_state_rsci_dout = {for_mux_127_nl , for_mux_126_nl , for_mux_125_nl ,
      for_mux_124_nl , for_mux_123_nl , for_mux_122_nl , for_mux_121_nl , for_mux_120_nl
      , for_mux_119_nl , for_mux_118_nl , for_mux_117_nl , for_mux_116_nl , for_mux_115_nl
      , for_mux_114_nl , for_mux_113_nl , for_mux_112_nl , for_mux_111_nl , for_mux_110_nl
      , for_mux_109_nl , for_mux_108_nl , for_mux_107_nl , for_mux_106_nl , for_mux_105_nl
      , for_mux_104_nl , for_mux_103_nl , for_mux_102_nl , for_mux_101_nl , for_mux_100_nl
      , for_mux_99_nl , for_mux_98_nl , for_mux_97_nl , for_mux_96_nl , for_mux_95_nl
      , for_mux_94_nl , for_mux_93_nl , for_mux_92_nl , for_mux_91_nl , for_mux_90_nl
      , for_mux_89_nl , for_mux_88_nl , for_mux_87_nl , for_mux_86_nl , for_mux_85_nl
      , for_mux_84_nl , for_mux_83_nl , for_mux_82_nl , for_mux_81_nl , for_mux_80_nl
      , for_mux_79_nl , for_mux_78_nl , for_mux_77_nl , for_mux_76_nl , for_mux_75_nl
      , for_mux_74_nl , for_mux_73_nl , for_mux_72_nl , for_mux_71_nl , for_mux_70_nl
      , for_mux_69_nl , for_mux_68_nl , for_mux_67_nl , for_mux_66_nl , for_mux_65_nl
      , for_mux_64_nl , for_mux_63_nl , for_mux_62_nl , for_mux_61_nl , for_mux_60_nl
      , for_mux_59_nl , for_mux_58_nl , for_mux_57_nl , for_mux_56_nl , for_mux_55_nl
      , for_mux_54_nl , for_mux_53_nl , for_mux_52_nl , for_mux_51_nl , for_mux_50_nl
      , for_mux_49_nl , for_mux_48_nl , for_mux_47_nl , for_mux_46_nl , for_mux_45_nl
      , for_mux_44_nl , for_mux_43_nl , for_mux_42_nl , for_mux_41_nl , for_mux_40_nl
      , for_mux_39_nl , for_mux_38_nl , for_mux_37_nl , for_mux_36_nl , for_mux_35_nl
      , for_mux_34_nl , for_mux_33_nl , for_mux_32_nl , for_mux_31_nl , for_mux_30_nl
      , for_mux_29_nl , for_mux_28_nl , for_mux_27_nl , for_mux_26_nl , for_mux_25_nl
      , for_mux_24_nl , for_mux_23_nl , for_mux_22_nl , for_mux_21_nl , for_mux_20_nl
      , for_mux_19_nl , for_mux_18_nl , for_mux_17_nl , for_mux_16_nl , for_mux_15_nl
      , for_mux_14_nl , for_mux_13_nl , for_mux_12_nl , for_mux_11_nl , for_mux_10_nl
      , for_mux_9_nl , for_mux_8_nl , for_mux_7_nl , for_mux_6_nl , for_mux_5_nl
      , for_mux_4_nl , for_mux_3_nl , for_mux_2_nl , for_mux_1_nl , for_mux_nl};
  wire  nl_MixColumns_core_core_fsm_inst_for_C_1_tr0;
  assign nl_MixColumns_core_core_fsm_inst_for_C_1_tr0 = i_2_0_sva_2[2];
  mgc_inout_prereg_en_v1 #(.rscid(32'sd1),
  .width(32'sd128)) state_rsci (
      .din(state_rsci_din),
      .ldout(nl_state_rsci_ldout),
      .dout(nl_state_rsci_dout[127:0]),
      .zin(state_rsc_zin),
      .lzout(state_rsc_lzout),
      .zout(state_rsc_zout)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) state_triosy_obj (
      .ld(state_triosy_obj_ld),
      .lz(state_triosy_lz)
    );
  MixColumns_core_core_fsm MixColumns_core_core_fsm_inst (
      .clk(clk),
      .rst_n(rst_n),
      .fsm_output(fsm_output),
      .for_C_1_tr0(nl_MixColumns_core_core_fsm_inst_for_C_1_tr0)
    );
  assign for_conc_35_cmx_7_sva_1 = (for_slc_state_8_7_0_4_ncse_sva_1[7]) ^ (for_slc_state_8_7_0_4_ncse_sva_1[6])
      ^ (t_sva_1[6]) ^ (Tmp_sva_1[7]);
  assign for_conc_35_cmx_6_sva_1 = (for_slc_state_8_7_0_4_ncse_sva_1[6]) ^ (for_slc_state_8_7_0_4_ncse_sva_1[5])
      ^ (t_sva_1[5]) ^ (Tmp_sva_1[6]);
  assign for_conc_35_cmx_5_sva_1 = (for_slc_state_8_7_0_4_ncse_sva_1[5]) ^ (for_slc_state_8_7_0_4_ncse_sva_1[4])
      ^ (t_sva_1[4]) ^ (Tmp_sva_1[5]);
  assign for_conc_32_cmx_2_sva_1 = (t_sva_1[2]) ^ (t_sva_1[1]) ^ (for_slc_state_8_7_0_2_cse_sva_1[1])
      ^ (Tmp_sva_1[2]);
  assign for_conc_35_cmx_2_sva_1 = (for_slc_state_8_7_0_4_ncse_sva_1[2]) ^ (for_slc_state_8_7_0_4_ncse_sva_1[1])
      ^ (t_sva_1[1]) ^ (Tmp_sva_1[2]);
  assign for_conc_32_cmx_5_sva_1 = (t_sva_1[5]) ^ (t_sva_1[4]) ^ (for_slc_state_8_7_0_2_cse_sva_1[4])
      ^ (Tmp_sva_1[5]);
  assign for_conc_32_cmx_6_sva_1 = (t_sva_1[6]) ^ (t_sva_1[5]) ^ (for_slc_state_8_7_0_2_cse_sva_1[5])
      ^ (Tmp_sva_1[6]);
  assign for_conc_32_cmx_7_sva_1 = (t_sva_1[7]) ^ (t_sva_1[6]) ^ (for_slc_state_8_7_0_2_cse_sva_1[6])
      ^ (Tmp_sva_1[7]);
  assign for_conc_34_cmx_7_sva_1 = (for_slc_state_8_7_0_3_ncse_sva_1[7]) ^ (for_slc_state_8_7_0_3_ncse_sva_1[6])
      ^ (for_slc_state_8_7_0_4_ncse_sva_1[6]) ^ (Tmp_sva_1[7]);
  assign for_conc_34_cmx_6_sva_1 = (for_slc_state_8_7_0_3_ncse_sva_1[6]) ^ (for_slc_state_8_7_0_3_ncse_sva_1[5])
      ^ (for_slc_state_8_7_0_4_ncse_sva_1[5]) ^ (Tmp_sva_1[6]);
  assign for_conc_34_cmx_5_sva_1 = (for_slc_state_8_7_0_3_ncse_sva_1[5]) ^ (for_slc_state_8_7_0_3_ncse_sva_1[4])
      ^ (for_slc_state_8_7_0_4_ncse_sva_1[4]) ^ (Tmp_sva_1[5]);
  assign for_conc_33_cmx_2_sva_1 = (for_slc_state_8_7_0_2_cse_sva_1[2]) ^ (for_slc_state_8_7_0_2_cse_sva_1[1])
      ^ (for_slc_state_8_7_0_3_ncse_sva_1[1]) ^ (Tmp_sva_1[2]);
  assign for_conc_34_cmx_2_sva_1 = (for_slc_state_8_7_0_3_ncse_sva_1[2]) ^ (for_slc_state_8_7_0_3_ncse_sva_1[1])
      ^ (for_slc_state_8_7_0_4_ncse_sva_1[1]) ^ (Tmp_sva_1[2]);
  assign for_conc_33_cmx_5_sva_1 = (for_slc_state_8_7_0_2_cse_sva_1[5]) ^ (for_slc_state_8_7_0_2_cse_sva_1[4])
      ^ (for_slc_state_8_7_0_3_ncse_sva_1[4]) ^ (Tmp_sva_1[5]);
  assign for_conc_33_cmx_6_sva_1 = (for_slc_state_8_7_0_2_cse_sva_1[6]) ^ (for_slc_state_8_7_0_2_cse_sva_1[5])
      ^ (for_slc_state_8_7_0_3_ncse_sva_1[5]) ^ (Tmp_sva_1[6]);
  assign for_conc_33_cmx_7_sva_1 = (for_slc_state_8_7_0_2_cse_sva_1[7]) ^ (for_slc_state_8_7_0_2_cse_sva_1[6])
      ^ (for_slc_state_8_7_0_3_ncse_sva_1[6]) ^ (Tmp_sva_1[7]);
  assign for_slc_state_8_7_0_4_ncse_sva_1 = MUX_v_8_4_2((state_rsci_din[31:24]),
      (state_rsci_din[63:56]), (state_rsci_din[95:88]), (state_rsci_din[127:120]),
      i_2_0_sva_1_0);
  assign t_sva_1 = MUX_v_8_4_2((state_rsci_din[7:0]), (state_rsci_din[39:32]), (state_rsci_din[71:64]),
      (state_rsci_din[103:96]), i_2_0_sva_1_0);
  assign Tmp_sva_1 = t_sva_1 ^ for_slc_state_8_7_0_2_cse_sva_1 ^ for_slc_state_8_7_0_3_ncse_sva_1
      ^ for_slc_state_8_7_0_4_ncse_sva_1;
  assign for_slc_state_8_7_0_3_ncse_sva_1 = MUX_v_8_4_2((state_rsci_din[23:16]),
      (state_rsci_din[55:48]), (state_rsci_din[87:80]), (state_rsci_din[119:112]),
      i_2_0_sva_1_0);
  assign for_slc_state_8_7_0_2_cse_sva_1 = MUX_v_8_4_2((state_rsci_din[15:8]), (state_rsci_din[47:40]),
      (state_rsci_din[79:72]), (state_rsci_din[111:104]), i_2_0_sva_1_0);
  assign nl_i_2_0_sva_2 = conv_u2u_2_3(i_2_0_sva_1_0) + 3'b001;
  assign i_2_0_sva_2 = nl_i_2_0_sva_2[2:0];
  assign and_dcpl = ~((i_2_0_sva_1_0!=2'b00));
  assign or_dcpl_1 = (i_2_0_sva_1_0!=2'b01);
  assign or_dcpl_2 = (i_2_0_sva_1_0!=2'b10);
  assign or_dcpl_3 = ~((i_2_0_sva_1_0==2'b11));
  assign for_conc_32_cmx_0_sva_1 = (t_sva_1[0]) ^ (t_sva_1[7]) ^ (for_slc_state_8_7_0_2_cse_sva_1[7])
      ^ (Tmp_sva_1[0]);
  assign xor_cse = (Tmp_sva_1[1]) ^ (t_sva_1[0]) ^ (t_sva_1[7]);
  assign for_conc_32_cmx_1_sva_1 = (t_sva_1[1]) ^ (for_slc_state_8_7_0_2_cse_sva_1[0])
      ^ (for_slc_state_8_7_0_2_cse_sva_1[7]) ^ xor_cse;
  assign xor_cse_1 = (for_slc_state_8_7_0_4_ncse_sva_1[7]) ^ (t_sva_1[7]) ^ (for_slc_state_8_7_0_4_ncse_sva_1[3]);
  assign for_conc_35_cmx_4_sva_1 = (t_sva_1[3]) ^ (for_slc_state_8_7_0_4_ncse_sva_1[4])
      ^ (Tmp_sva_1[4]) ^ xor_cse_1;
  assign xor_cse_2 = (for_slc_state_8_7_0_2_cse_sva_1[7]) ^ (t_sva_1[7]) ^ (t_sva_1[3]);
  assign for_conc_32_cmx_3_sva_1 = (t_sva_1[2]) ^ (for_slc_state_8_7_0_2_cse_sva_1[2])
      ^ (Tmp_sva_1[3]) ^ xor_cse_2;
  assign for_conc_35_cmx_3_sva_1 = (for_slc_state_8_7_0_4_ncse_sva_1[2]) ^ (t_sva_1[2])
      ^ (Tmp_sva_1[3]) ^ xor_cse_1;
  assign for_conc_32_cmx_4_sva_1 = (for_slc_state_8_7_0_2_cse_sva_1[3]) ^ (t_sva_1[4])
      ^ (Tmp_sva_1[4]) ^ xor_cse_2;
  assign for_conc_35_cmx_1_sva_1 = (for_slc_state_8_7_0_4_ncse_sva_1[1]) ^ (for_slc_state_8_7_0_4_ncse_sva_1[0])
      ^ (for_slc_state_8_7_0_4_ncse_sva_1[7]) ^ xor_cse;
  assign for_conc_35_cmx_0_sva_1 = (for_slc_state_8_7_0_4_ncse_sva_1[0]) ^ (for_slc_state_8_7_0_4_ncse_sva_1[7])
      ^ (t_sva_1[7]) ^ (Tmp_sva_1[0]);
  assign for_conc_33_cmx_0_sva_1 = (for_slc_state_8_7_0_2_cse_sva_1[0]) ^ (for_slc_state_8_7_0_2_cse_sva_1[7])
      ^ (for_slc_state_8_7_0_3_ncse_sva_1[7]) ^ (Tmp_sva_1[0]);
  assign xor_cse_3 = (for_slc_state_8_7_0_3_ncse_sva_1[7]) ^ (for_slc_state_8_7_0_3_ncse_sva_1[0])
      ^ (Tmp_sva_1[1]);
  assign for_conc_33_cmx_1_sva_1 = (for_slc_state_8_7_0_2_cse_sva_1[1]) ^ (for_slc_state_8_7_0_2_cse_sva_1[0])
      ^ (for_slc_state_8_7_0_2_cse_sva_1[7]) ^ xor_cse_3;
  assign xor_cse_4 = (for_slc_state_8_7_0_4_ncse_sva_1[7]) ^ (for_slc_state_8_7_0_3_ncse_sva_1[7])
      ^ (for_slc_state_8_7_0_3_ncse_sva_1[3]);
  assign for_conc_34_cmx_4_sva_1 = (for_slc_state_8_7_0_4_ncse_sva_1[3]) ^ (for_slc_state_8_7_0_3_ncse_sva_1[4])
      ^ (Tmp_sva_1[4]) ^ xor_cse_4;
  assign xor_cse_5 = (for_slc_state_8_7_0_3_ncse_sva_1[7]) ^ (for_slc_state_8_7_0_2_cse_sva_1[7])
      ^ (for_slc_state_8_7_0_2_cse_sva_1[3]);
  assign for_conc_33_cmx_3_sva_1 = (for_slc_state_8_7_0_2_cse_sva_1[2]) ^ (for_slc_state_8_7_0_3_ncse_sva_1[2])
      ^ (Tmp_sva_1[3]) ^ xor_cse_5;
  assign for_conc_34_cmx_3_sva_1 = (for_slc_state_8_7_0_3_ncse_sva_1[2]) ^ (for_slc_state_8_7_0_4_ncse_sva_1[2])
      ^ (Tmp_sva_1[3]) ^ xor_cse_4;
  assign for_conc_33_cmx_4_sva_1 = (for_slc_state_8_7_0_3_ncse_sva_1[3]) ^ (for_slc_state_8_7_0_2_cse_sva_1[4])
      ^ (Tmp_sva_1[4]) ^ xor_cse_5;
  assign for_conc_34_cmx_1_sva_1 = (for_slc_state_8_7_0_3_ncse_sva_1[1]) ^ (for_slc_state_8_7_0_4_ncse_sva_1[0])
      ^ (for_slc_state_8_7_0_4_ncse_sva_1[7]) ^ xor_cse_3;
  assign for_conc_34_cmx_0_sva_1 = (for_slc_state_8_7_0_3_ncse_sva_1[0]) ^ (for_slc_state_8_7_0_3_ncse_sva_1[7])
      ^ (for_slc_state_8_7_0_4_ncse_sva_1[7]) ^ (Tmp_sva_1[0]);
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      i_2_0_sva_1_0 <= 2'b00;
    end
    else if ( (fsm_output[0]) | (fsm_output[2]) ) begin
      i_2_0_sva_1_0 <= MUX_v_2_2_2(2'b00, (i_2_0_sva_2[1:0]), i_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      state_triosy_obj_ld <= 1'b0;
    end
    else begin
      state_triosy_obj_ld <= (i_2_0_sva_2[2]) & (fsm_output[2]);
    end
  end
  assign i_not_1_nl = ~ (fsm_output[0]);

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_4_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [1:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_8_4_2 = result;
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MixColumns
// ------------------------------------------------------------------


module MixColumns (
  clk, rst_n, state_rsc_zout, state_rsc_lzout, state_rsc_zin, state_triosy_lz
);
  input clk;
  input rst_n;
  output [127:0] state_rsc_zout;
  output state_rsc_lzout;
  input [127:0] state_rsc_zin;
  output state_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  MixColumns_core MixColumns_core_inst (
      .clk(clk),
      .rst_n(rst_n),
      .state_rsc_zout(state_rsc_zout),
      .state_rsc_lzout(state_rsc_lzout),
      .state_rsc_zin(state_rsc_zin),
      .state_triosy_lz(state_triosy_lz)
    );
endmodule



