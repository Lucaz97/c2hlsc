
//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_inout_prereg_en_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2019 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_inout_prereg_en_v1 (din, ldout, dout, zin, lzout, zout);

    parameter integer rscid = 1;
    parameter integer width = 8;

    output [width-1:0] din;
    input              ldout;
    input  [width-1:0] dout;
    input  [width-1:0] zin;
    output             lzout;
    output [width-1:0] zout;

    wire   [width-1:0] din;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzout = ldout;
    assign din = zin;
    assign zout = dout;

endmodule



//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   lc4976@hansolo.poly.edu
//  Generated date: Tue Apr  9 22:15:36 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    quickSort_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module quickSort_core_core_fsm (
  clk, rst_n, fsm_output, while_C_0_tr0, partition_while_while_C_0_tr0, partition_while_while_1_C_0_tr0,
      partition_while_C_1_tr0, while_C_3_tr0
);
  input clk;
  input rst_n;
  output [11:0] fsm_output;
  reg [11:0] fsm_output;
  input while_C_0_tr0;
  input partition_while_while_C_0_tr0;
  input partition_while_while_1_C_0_tr0;
  input partition_while_C_1_tr0;
  input while_C_3_tr0;


  // FSM State Type Declaration for quickSort_core_core_fsm_1
  parameter
    main_C_0 = 4'd0,
    while_C_0 = 4'd1,
    partition_while_while_C_0 = 4'd2,
    partition_while_while_C_1 = 4'd3,
    partition_while_while_1_C_0 = 4'd4,
    partition_while_while_1_C_1 = 4'd5,
    partition_while_C_0 = 4'd6,
    partition_while_C_1 = 4'd7,
    while_C_1 = 4'd8,
    while_C_2 = 4'd9,
    while_C_3 = 4'd10,
    main_C_1 = 4'd11;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : quickSort_core_core_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 12'b000000000010;
        if ( while_C_0_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = partition_while_while_C_0;
        end
      end
      partition_while_while_C_0 : begin
        fsm_output = 12'b000000000100;
        if ( partition_while_while_C_0_tr0 ) begin
          state_var_NS = partition_while_while_1_C_0;
        end
        else begin
          state_var_NS = partition_while_while_C_1;
        end
      end
      partition_while_while_C_1 : begin
        fsm_output = 12'b000000001000;
        state_var_NS = partition_while_while_C_0;
      end
      partition_while_while_1_C_0 : begin
        fsm_output = 12'b000000010000;
        if ( partition_while_while_1_C_0_tr0 ) begin
          state_var_NS = partition_while_C_0;
        end
        else begin
          state_var_NS = partition_while_while_1_C_1;
        end
      end
      partition_while_while_1_C_1 : begin
        fsm_output = 12'b000000100000;
        state_var_NS = partition_while_while_1_C_0;
      end
      partition_while_C_0 : begin
        fsm_output = 12'b000001000000;
        state_var_NS = partition_while_C_1;
      end
      partition_while_C_1 : begin
        fsm_output = 12'b000010000000;
        if ( partition_while_C_1_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = partition_while_while_C_0;
        end
      end
      while_C_1 : begin
        fsm_output = 12'b000100000000;
        state_var_NS = while_C_2;
      end
      while_C_2 : begin
        fsm_output = 12'b001000000000;
        state_var_NS = while_C_3;
      end
      while_C_3 : begin
        fsm_output = 12'b010000000000;
        if ( while_C_3_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 12'b100000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 12'b000000000001;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    quickSort_core
// ------------------------------------------------------------------


module quickSort_core (
  clk, rst_n, arr_rsc_zout, arr_rsc_lzout, arr_rsc_zin, arr_triosy_lz, low_rsc_dat,
      low_triosy_lz, high_rsc_dat, high_triosy_lz
);
  input clk;
  input rst_n;
  output [2047:0] arr_rsc_zout;
  output arr_rsc_lzout;
  input [2047:0] arr_rsc_zin;
  output arr_triosy_lz;
  input [31:0] low_rsc_dat;
  output low_triosy_lz;
  input [31:0] high_rsc_dat;
  output high_triosy_lz;


  // Interconnect Declarations
  wire [2047:0] arr_rsci_din;
  wire [31:0] low_rsci_idat;
  wire [31:0] high_rsci_idat;
  wire [11:0] fsm_output;
  wire [29:0] while_if_slc_while_if_while_if_acc_tmp;
  wire [30:0] nl_while_if_slc_while_if_while_if_acc_tmp;
  wire or_dcpl_1;
  wire and_dcpl;
  wire and_dcpl_73;
  wire or_tmp_613;
  reg exit_partition_while_sva;
  wire swap_1_equal_tmp_283;
  wire swap_1_equal_tmp_285;
  reg swap_1_equal_tmp_3;
  wire swap_1_equal_tmp_288;
  reg swap_1_equal_tmp_5;
  wire swap_1_equal_tmp_291;
  reg swap_1_equal_tmp_7;
  wire swap_1_equal_tmp_293;
  wire swap_1_equal_tmp_295;
  reg swap_1_equal_tmp_11;
  wire swap_1_equal_tmp_296;
  reg swap_1_equal_tmp_13;
  reg swap_1_equal_tmp_14;
  reg swap_1_equal_tmp_15;
  wire swap_1_equal_tmp_298;
  reg swap_1_equal_tmp_17;
  reg swap_1_equal_tmp_18;
  reg swap_1_equal_tmp_19;
  reg swap_1_equal_tmp_20;
  reg swap_1_equal_tmp_21;
  reg swap_1_equal_tmp_22;
  reg swap_1_equal_tmp_23;
  reg swap_1_equal_tmp_24;
  reg swap_1_equal_tmp_25;
  reg swap_1_equal_tmp_26;
  reg swap_1_equal_tmp_27;
  reg swap_1_equal_tmp_28;
  reg swap_1_equal_tmp_29;
  reg swap_1_equal_tmp_30;
  reg swap_1_equal_tmp_31;
  wire swap_1_equal_tmp_305;
  reg swap_1_equal_tmp_33;
  reg swap_1_equal_tmp_34;
  reg swap_1_equal_tmp_35;
  reg swap_1_equal_tmp_36;
  reg swap_1_equal_tmp_37;
  reg swap_1_equal_tmp_38;
  reg swap_1_equal_tmp_39;
  reg swap_1_equal_tmp_40;
  reg swap_1_equal_tmp_41;
  reg swap_1_equal_tmp_42;
  reg swap_1_equal_tmp_43;
  reg swap_1_equal_tmp_44;
  reg swap_1_equal_tmp_45;
  reg swap_1_equal_tmp_46;
  reg swap_1_equal_tmp_47;
  reg swap_1_equal_tmp_48;
  reg swap_1_equal_tmp_49;
  reg swap_1_equal_tmp_50;
  reg swap_1_equal_tmp_51;
  reg swap_1_equal_tmp_52;
  reg swap_1_equal_tmp_53;
  reg swap_1_equal_tmp_54;
  reg swap_1_equal_tmp_55;
  reg swap_1_equal_tmp_56;
  reg swap_1_equal_tmp_57;
  reg swap_1_equal_tmp_58;
  reg swap_1_equal_tmp_59;
  reg swap_1_equal_tmp_60;
  reg swap_1_equal_tmp_61;
  reg swap_1_equal_tmp_62;
  reg swap_1_equal_tmp_63;
  wire swap_1_equal_tmp_284;
  wire swap_1_equal_tmp_286;
  wire swap_1_equal_tmp_287;
  wire swap_1_equal_tmp_289;
  wire swap_1_equal_tmp_290;
  wire swap_1_equal_tmp_292;
  reg swap_1_equal_tmp_71;
  wire swap_1_equal_tmp_294;
  reg swap_1_equal_tmp_73;
  reg swap_1_equal_tmp_74;
  reg swap_1_equal_tmp_75;
  reg swap_1_equal_tmp_76;
  reg swap_1_equal_tmp_77;
  reg swap_1_equal_tmp_78;
  reg swap_1_equal_tmp_79;
  wire swap_1_equal_tmp_299;
  wire swap_1_equal_tmp_300;
  wire swap_1_equal_tmp_301;
  reg swap_1_equal_tmp_83;
  wire swap_1_equal_tmp_302;
  reg swap_1_equal_tmp_85;
  reg swap_1_equal_tmp_86;
  reg swap_1_equal_tmp_87;
  reg swap_1_equal_tmp_88;
  reg swap_1_equal_tmp_89;
  reg swap_1_equal_tmp_90;
  reg swap_1_equal_tmp_91;
  reg swap_1_equal_tmp_92;
  reg swap_1_equal_tmp_93;
  reg swap_1_equal_tmp_94;
  reg swap_1_equal_tmp_95;
  wire swap_1_equal_tmp_306;
  reg swap_1_equal_tmp_97;
  wire swap_1_equal_tmp_304;
  reg swap_1_equal_tmp_99;
  reg swap_1_equal_tmp_100;
  reg swap_1_equal_tmp_101;
  reg swap_1_equal_tmp_102;
  reg swap_1_equal_tmp_103;
  wire swap_1_equal_tmp_303;
  reg swap_1_equal_tmp_105;
  reg swap_1_equal_tmp_106;
  reg swap_1_equal_tmp_107;
  reg swap_1_equal_tmp_108;
  reg swap_1_equal_tmp_109;
  reg swap_1_equal_tmp_110;
  reg swap_1_equal_tmp_111;
  wire swap_1_equal_tmp_297;
  reg swap_1_equal_tmp_113;
  reg swap_1_equal_tmp_114;
  reg swap_1_equal_tmp_115;
  reg swap_1_equal_tmp_116;
  reg swap_1_equal_tmp_117;
  reg swap_1_equal_tmp_118;
  reg swap_1_equal_tmp_119;
  reg swap_1_equal_tmp_120;
  reg swap_1_equal_tmp_121;
  reg swap_1_equal_tmp_122;
  reg swap_1_equal_tmp_123;
  reg swap_1_equal_tmp_124;
  reg swap_1_equal_tmp_125;
  reg swap_1_equal_tmp_126;
  reg swap_1_equal_tmp_127;
  reg swap_1_nor_101_itm;
  reg swap_1_nor_94_itm;
  reg swap_1_nor_88_itm;
  reg swap_1_nor_86_itm;
  reg swap_1_nor_75_itm;
  reg swap_1_nor_73_itm;
  reg swap_1_nor_72_itm;
  reg swap_1_nor_71_itm;
  reg swap_1_nor_63_itm;
  reg swap_1_nor_61_itm;
  reg swap_1_nor_60_itm;
  reg swap_1_nor_59_itm;
  reg swap_1_nor_58_itm;
  reg swap_1_nor_57_itm;
  reg swap_1_nor_56_itm;
  reg swap_1_nor_30_itm;
  reg swap_1_nor_15_itm;
  reg swap_1_nor_11_itm;
  reg swap_1_nor_8_itm;
  reg swap_1_nor_7_itm;
  reg swap_1_nor_5_itm;
  reg swap_1_nor_3_itm;
  reg swap_1_nor_1_itm;
  reg swap_1_nor_itm;
  wire swap_equal_tmp_178;
  wire swap_equal_tmp_181;
  wire swap_equal_tmp_184;
  wire swap_equal_tmp_187;
  wire swap_equal_tmp_190;
  wire swap_equal_tmp_193;
  wire swap_equal_tmp_196;
  wire swap_equal_tmp_198;
  wire swap_equal_tmp_201;
  wire swap_equal_tmp_203;
  wire swap_equal_tmp_205;
  wire swap_equal_tmp_207;
  wire swap_equal_tmp_209;
  wire swap_equal_tmp_211;
  wire swap_equal_tmp_214;
  wire swap_equal_tmp_216;
  wire swap_equal_tmp_219;
  wire swap_equal_tmp_222;
  wire swap_equal_tmp_225;
  wire swap_equal_tmp_227;
  wire swap_equal_tmp_230;
  wire swap_equal_tmp_232;
  wire swap_equal_tmp_235;
  wire swap_equal_tmp_237;
  wire swap_equal_tmp_239;
  wire swap_equal_tmp_241;
  wire swap_equal_tmp_243;
  wire swap_equal_tmp_245;
  wire swap_equal_tmp_248;
  wire swap_equal_tmp_250;
  wire swap_equal_tmp_253;
  wire swap_equal_tmp_251;
  wire swap_equal_tmp_249;
  wire swap_equal_tmp_246;
  wire swap_equal_tmp_244;
  wire swap_equal_tmp_242;
  wire swap_equal_tmp_240;
  wire swap_equal_tmp_238;
  wire swap_equal_tmp_236;
  wire swap_equal_tmp_233;
  wire swap_equal_tmp_231;
  wire swap_equal_tmp_229;
  wire swap_equal_tmp_226;
  wire swap_equal_tmp_224;
  wire swap_equal_tmp_221;
  wire swap_equal_tmp_218;
  wire swap_equal_tmp_215;
  wire swap_equal_tmp_212;
  wire swap_equal_tmp_210;
  wire swap_equal_tmp_208;
  wire swap_equal_tmp_206;
  wire swap_equal_tmp_204;
  wire swap_equal_tmp_202;
  wire swap_equal_tmp_200;
  wire swap_equal_tmp_197;
  wire swap_equal_tmp_195;
  wire swap_equal_tmp_192;
  wire swap_equal_tmp_189;
  wire swap_equal_tmp_186;
  wire swap_equal_tmp_183;
  wire swap_equal_tmp_180;
  wire swap_equal_tmp_177;
  wire swap_equal_tmp_176;
  wire swap_equal_tmp_179;
  wire swap_equal_tmp_182;
  wire swap_equal_tmp_185;
  wire swap_equal_tmp_188;
  wire swap_equal_tmp_191;
  wire swap_equal_tmp_194;
  wire swap_equal_tmp_136;
  wire swap_equal_tmp_199;
  wire swap_equal_tmp_139;
  wire swap_equal_tmp_141;
  wire swap_equal_tmp_143;
  wire swap_equal_tmp_145;
  wire swap_equal_tmp_147;
  wire swap_equal_tmp_149;
  wire swap_equal_tmp_150;
  wire swap_equal_tmp_217;
  wire swap_equal_tmp_220;
  wire swap_equal_tmp_223;
  wire swap_equal_tmp_155;
  wire swap_equal_tmp_228;
  wire swap_equal_tmp_158;
  wire swap_equal_tmp_160;
  wire swap_equal_tmp_161;
  wire swap_equal_tmp_163;
  wire swap_equal_tmp_165;
  wire swap_equal_tmp_167;
  wire swap_equal_tmp_169;
  wire swap_equal_tmp_171;
  wire swap_equal_tmp_172;
  wire swap_equal_tmp_174;
  wire swap_equal_tmp_175;
  wire swap_equal_tmp_252;
  wire swap_equal_tmp_173;
  wire swap_equal_tmp_247;
  wire swap_equal_tmp_170;
  wire swap_equal_tmp_168;
  wire swap_equal_tmp_166;
  wire swap_equal_tmp_164;
  wire swap_equal_tmp_162;
  wire swap_equal_tmp_234;
  wire swap_equal_tmp_159;
  wire swap_equal_tmp_157;
  wire swap_equal_tmp_156;
  wire swap_equal_tmp_154;
  wire swap_equal_tmp_153;
  wire swap_equal_tmp_152;
  wire swap_equal_tmp_151;
  wire swap_equal_tmp_213;
  wire swap_equal_tmp_148;
  wire swap_equal_tmp_146;
  wire swap_equal_tmp_144;
  wire swap_equal_tmp_142;
  wire swap_equal_tmp_140;
  wire swap_equal_tmp_138;
  wire swap_equal_tmp_137;
  wire swap_equal_tmp_135;
  wire swap_equal_tmp_134;
  wire swap_equal_tmp_133;
  wire swap_equal_tmp_132;
  wire swap_equal_tmp_131;
  wire swap_equal_tmp_130;
  wire swap_equal_tmp_129;
  wire swap_equal_tmp_128;
  wire swap_1_nor_101_itm_1;
  wire swap_1_nor_94_itm_2;
  wire swap_1_nor_88_itm_2;
  wire swap_1_nor_86_itm_2;
  wire swap_1_nor_75_itm_2;
  wire swap_1_nor_73_itm_2;
  wire swap_1_nor_72_itm_2;
  wire swap_1_nor_71_itm_2;
  wire swap_1_nor_63_itm_2;
  wire swap_1_nor_61_itm_2;
  wire swap_1_nor_60_itm_2;
  wire swap_1_nor_59_itm_2;
  wire swap_1_nor_58_itm_1;
  wire swap_1_nor_57_itm_1;
  wire swap_1_nor_56_itm_1;
  reg [31:0] partition_j_lpi_4;
  reg [31:0] partition_i_lpi_4;
  reg [31:0] stack_0_1_sva;
  reg [31:0] stack_2_1_sva;
  reg [31:0] stack_4_1_sva;
  reg [31:0] stack_6_1_sva;
  reg [31:0] stack_8_1_sva;
  reg [31:0] stack_10_1_sva;
  reg [31:0] stack_12_1_sva;
  reg [31:0] stack_14_1_sva;
  reg [31:0] stack_16_1_sva;
  reg [31:0] stack_18_1_sva;
  reg [31:0] stack_20_1_sva;
  reg [31:0] stack_22_1_sva;
  reg [31:0] stack_24_1_sva;
  reg [31:0] stack_26_1_sva;
  reg [31:0] stack_28_1_sva;
  reg [31:0] stack_30_1_sva;
  reg [31:0] stack_32_1_sva;
  reg [31:0] stack_34_1_sva;
  reg [31:0] stack_36_1_sva;
  reg [31:0] stack_38_1_sva;
  reg [31:0] stack_40_1_sva;
  reg [31:0] stack_42_1_sva;
  reg [31:0] stack_44_1_sva;
  reg [31:0] stack_46_1_sva;
  reg [31:0] stack_48_1_sva;
  reg [31:0] stack_50_1_sva;
  reg [31:0] stack_52_1_sva;
  reg [31:0] stack_54_1_sva;
  reg [31:0] stack_56_1_sva;
  reg [31:0] stack_58_1_sva;
  reg [31:0] stack_60_1_sva;
  reg [31:0] stack_62_1_sva;
  reg [31:0] stack_64_1_sva;
  reg [31:0] stack_66_1_sva;
  reg [31:0] stack_68_1_sva;
  reg [31:0] stack_70_1_sva;
  reg [31:0] stack_72_1_sva;
  reg [31:0] stack_74_1_sva;
  reg [31:0] stack_76_1_sva;
  reg [31:0] stack_78_1_sva;
  reg [31:0] stack_80_1_sva;
  reg [31:0] stack_82_1_sva;
  reg [31:0] stack_84_1_sva;
  reg [31:0] stack_86_1_sva;
  reg [31:0] stack_88_1_sva;
  reg [31:0] stack_90_1_sva;
  reg [31:0] stack_92_1_sva;
  reg [31:0] stack_94_1_sva;
  reg [31:0] stack_96_1_sva;
  reg [31:0] stack_98_1_sva;
  reg [31:0] stack_100_1_sva;
  reg [31:0] stack_102_1_sva;
  reg [31:0] stack_104_1_sva;
  reg [31:0] stack_106_1_sva;
  reg [31:0] stack_108_1_sva;
  reg [31:0] stack_110_1_sva;
  reg [31:0] stack_112_1_sva;
  reg [31:0] stack_114_1_sva;
  reg [31:0] stack_116_1_sva;
  reg [31:0] stack_118_1_sva;
  reg [31:0] stack_120_1_sva;
  reg [31:0] stack_122_1_sva;
  reg [31:0] stack_124_1_sva;
  reg [31:0] stack_126_1_sva;
  reg [31:0] stack_1_1_sva;
  reg [31:0] stack_3_1_sva;
  reg [31:0] stack_5_1_sva;
  reg [31:0] stack_7_1_sva;
  reg [31:0] stack_9_1_sva;
  reg [31:0] stack_11_1_sva;
  reg [31:0] stack_13_1_sva;
  reg [31:0] stack_15_1_sva;
  reg [31:0] stack_17_1_sva;
  reg [31:0] stack_19_1_sva;
  reg [31:0] stack_21_1_sva;
  reg [31:0] stack_23_1_sva;
  reg [31:0] stack_25_1_sva;
  reg [31:0] stack_27_1_sva;
  reg [31:0] stack_29_1_sva;
  reg [31:0] stack_31_1_sva;
  reg [31:0] stack_33_1_sva;
  reg [31:0] stack_35_1_sva;
  reg [31:0] stack_37_1_sva;
  reg [31:0] stack_39_1_sva;
  reg [31:0] stack_41_1_sva;
  reg [31:0] stack_43_1_sva;
  reg [31:0] stack_45_1_sva;
  reg [31:0] stack_47_1_sva;
  reg [31:0] stack_49_1_sva;
  reg [31:0] stack_51_1_sva;
  reg [31:0] stack_53_1_sva;
  reg [31:0] stack_55_1_sva;
  reg [31:0] stack_57_1_sva;
  reg [31:0] stack_59_1_sva;
  reg [31:0] stack_61_1_sva;
  reg [31:0] stack_63_1_sva;
  reg [31:0] stack_65_1_sva;
  reg [31:0] stack_67_1_sva;
  reg [31:0] stack_69_1_sva;
  reg [31:0] stack_71_1_sva;
  reg [31:0] stack_73_1_sva;
  reg [31:0] stack_75_1_sva;
  reg [31:0] stack_77_1_sva;
  reg [31:0] stack_79_1_sva;
  reg [31:0] stack_81_1_sva;
  reg [31:0] stack_83_1_sva;
  reg [31:0] stack_85_1_sva;
  reg [31:0] stack_87_1_sva;
  reg [31:0] stack_89_1_sva;
  reg [31:0] stack_91_1_sva;
  reg [31:0] stack_93_1_sva;
  reg [31:0] stack_95_1_sva;
  reg [31:0] stack_97_1_sva;
  reg [31:0] stack_99_1_sva;
  reg [31:0] stack_101_1_sva;
  reg [31:0] stack_103_1_sva;
  reg [31:0] stack_105_1_sva;
  reg [31:0] stack_107_1_sva;
  reg [31:0] stack_109_1_sva;
  reg [31:0] stack_111_1_sva;
  reg [31:0] stack_113_1_sva;
  reg [31:0] stack_115_1_sva;
  reg [31:0] stack_117_1_sva;
  reg [31:0] stack_119_1_sva;
  reg [31:0] stack_121_1_sva;
  reg [31:0] stack_123_1_sva;
  reg [31:0] stack_125_1_sva;
  reg [31:0] stack_127_1_sva;
  reg while_acc_3_cse_32;
  wire while_if_and_stg_4_30_sva_1;
  wire while_if_and_stg_4_1_sva_1;
  wire while_if_and_stg_4_29_sva_1;
  wire while_if_and_stg_4_2_sva_1;
  wire while_if_and_stg_4_28_sva_1;
  wire while_if_and_stg_4_3_sva_1;
  wire while_if_and_stg_4_27_sva_1;
  wire while_if_and_stg_4_4_sva_1;
  wire while_if_and_stg_4_26_sva_1;
  wire while_if_and_stg_4_5_sva_1;
  wire while_if_and_stg_4_25_sva_1;
  wire while_if_and_stg_4_6_sva_1;
  wire while_if_and_stg_4_24_sva_1;
  wire while_if_and_stg_4_7_sva_1;
  wire while_if_and_stg_4_23_sva_1;
  wire while_if_and_stg_4_8_sva_1;
  wire while_if_and_stg_4_22_sva_1;
  wire while_if_and_stg_4_9_sva_1;
  wire while_if_and_stg_4_21_sva_1;
  wire while_if_and_stg_4_10_sva_1;
  wire while_if_and_stg_4_20_sva_1;
  wire while_if_and_stg_4_11_sva_1;
  wire while_if_and_stg_4_19_sva_1;
  wire while_if_and_stg_4_12_sva_1;
  wire while_if_and_stg_4_18_sva_1;
  wire while_if_and_stg_4_13_sva_1;
  wire while_if_and_stg_4_17_sva_1;
  wire while_if_and_stg_4_14_sva_1;
  wire while_if_and_stg_4_16_sva_1;
  wire while_if_and_stg_4_15_sva_1;
  wire while_if_and_stg_3_1_sva_1;
  wire while_if_and_stg_3_2_sva_1;
  wire while_if_and_stg_3_3_sva_1;
  wire while_if_and_stg_3_4_sva_1;
  wire while_if_and_stg_3_5_sva_1;
  wire while_if_and_stg_3_6_sva_1;
  wire while_if_and_stg_3_7_sva_1;
  wire while_if_and_stg_3_8_sva_1;
  wire while_if_and_stg_3_9_sva_1;
  wire while_if_and_stg_3_10_sva_1;
  wire while_if_and_stg_3_11_sva_1;
  wire while_if_and_stg_3_12_sva_1;
  wire while_if_and_stg_3_13_sva_1;
  wire while_if_and_stg_3_14_sva_1;
  wire while_if_and_stg_2_1_sva_1;
  wire while_if_and_stg_2_2_sva_1;
  wire while_if_and_stg_2_3_sva_1;
  wire while_if_and_stg_2_4_sva_1;
  wire while_if_and_stg_2_5_sva_1;
  wire while_if_and_stg_2_6_sva_1;
  wire while_if_and_stg_1_1_sva_1;
  wire while_if_and_stg_1_2_sva_1;
  wire while_if_and_369_tmp_sva_1;
  wire while_if_and_122_tmp_sva_1;
  wire while_if_and_stg_4_31_sva_1;
  wire while_if_and_stg_4_0_sva_1;
  wire while_if_and_stg_3_0_sva_1;
  wire while_if_and_stg_2_0_sva_1;
  wire while_if_and_stg_1_0_sva_1;
  wire while_if_and_stg_3_15_sva_1;
  wire while_if_and_stg_2_7_sva_1;
  wire while_if_and_stg_1_3_sva_1;
  reg [30:0] top_1_31_1_sva_1;
  reg while_if_slc_while_if_while_if_acc_1_psp_sva_5;
  wire [31:0] partition_while_while_1_mux_2;
  reg [31:0] low_sva;
  reg [31:0] high_sva;
  reg reg_high_triosy_obj_ld_cse;
  reg [1:0] partition_pivot_sva_31_30;
  reg [29:0] partition_pivot_sva_29_0;
  wire swap_or_64_tmp_1;
  wire swap_or_tmp_1;
  wire swap_1_or_tmp_1;
  wire swap_1_or_64_tmp_1;
  wire [31:0] z_out;
  wire or_tmp_637;
  wire [32:0] z_out_1;
  wire [31:0] low_sva_1;
  wire [31:0] high_sva_1;
  wire while_asn_523;
  wire while_asn_525;
  wire while_asn_529;
  wire while_asn_533;
  wire while_asn_537;
  wire while_asn_541;
  wire while_asn_545;
  wire while_asn_549;
  wire while_asn_553;
  wire while_asn_557;
  wire while_asn_561;
  wire while_asn_565;
  wire while_asn_569;
  wire while_asn_573;
  wire while_asn_577;
  wire while_asn_581;
  wire while_asn_585;
  wire while_asn_589;
  wire while_asn_593;
  wire while_asn_597;
  wire while_asn_601;
  wire while_asn_605;
  wire while_asn_609;
  wire while_asn_613;
  wire while_asn_617;
  wire while_asn_621;
  wire while_asn_625;
  wire while_asn_629;
  wire while_asn_633;
  wire while_asn_637;
  wire while_asn_641;
  wire while_asn_645;
  wire while_asn_649;
  wire while_asn_653;
  wire while_asn_657;
  wire while_asn_661;
  wire while_asn_665;
  wire while_asn_669;
  wire while_asn_673;
  wire while_asn_677;
  wire while_asn_681;
  wire while_asn_685;
  wire while_asn_689;
  wire while_asn_693;
  wire while_asn_697;
  wire while_asn_701;
  wire while_asn_705;
  wire while_asn_709;
  wire while_asn_713;
  wire while_asn_717;
  wire while_asn_721;
  wire while_asn_725;
  wire while_asn_729;
  wire while_asn_733;
  wire while_asn_737;
  wire while_asn_741;
  wire while_asn_745;
  wire while_asn_749;
  wire while_asn_753;
  wire while_asn_757;
  wire while_asn_761;
  wire while_asn_765;
  wire while_asn_769;
  wire while_asn_773;
  wire while_and_1_rgt;
  wire while_or_193_ssc;
  wire while_or_191_ssc;
  wire stack_and_1_cse;
  wire stack_and_2_cse;
  wire stack_and_3_cse;
  wire stack_and_4_cse;
  wire stack_and_5_cse;
  wire stack_and_6_cse;
  wire stack_and_7_cse;
  wire stack_and_8_cse;
  wire stack_and_9_cse;
  wire stack_and_10_cse;
  wire stack_and_11_cse;
  wire stack_and_12_cse;
  wire stack_and_13_cse;
  wire stack_and_14_cse;
  wire stack_and_15_cse;
  wire stack_and_16_cse;
  wire stack_and_17_cse;
  wire stack_and_18_cse;
  wire stack_and_19_cse;
  wire stack_and_20_cse;
  wire stack_and_21_cse;
  wire stack_and_22_cse;
  wire stack_and_23_cse;
  wire stack_and_24_cse;
  wire stack_and_25_cse;
  wire stack_and_26_cse;
  wire stack_and_27_cse;
  wire stack_and_28_cse;
  wire stack_and_29_cse;
  wire stack_and_30_cse;
  wire stack_and_31_cse;
  wire stack_and_32_cse;
  wire stack_and_33_cse;
  wire stack_and_34_cse;
  wire stack_and_35_cse;
  wire stack_and_36_cse;
  wire stack_and_37_cse;
  wire stack_and_38_cse;
  wire stack_and_39_cse;
  wire stack_and_40_cse;
  wire stack_and_41_cse;
  wire stack_and_42_cse;
  wire stack_and_43_cse;
  wire stack_and_44_cse;
  wire stack_and_45_cse;
  wire stack_and_46_cse;
  wire stack_and_47_cse;
  wire stack_and_48_cse;
  wire stack_and_49_cse;
  wire stack_and_50_cse;
  wire stack_and_51_cse;
  wire stack_and_52_cse;
  wire stack_and_53_cse;
  wire stack_and_54_cse;
  wire stack_and_55_cse;
  wire stack_and_56_cse;
  wire stack_and_57_cse;
  wire stack_and_58_cse;
  wire stack_and_59_cse;
  wire stack_and_60_cse;
  wire stack_and_61_cse;
  wire stack_and_62_cse;
  wire stack_and_63_cse;
  wire nand_87_cse;
  wire while_acc_3_itm_32_1;
  wire z_out_2_32;

  wire and_1186_nl;
  wire and_1187_nl;
  wire and_1188_nl;
  wire and_1189_nl;
  wire[29:0] and_1160_nl;
  wire[29:0] mux_nl;
  wire or_779_nl;
  wire or_747_nl;
  wire swap_1_nor_30_nl;
  wire swap_1_nor_15_nl;
  wire swap_1_nor_11_nl;
  wire swap_1_nor_5_nl;
  wire swap_1_nor_3_nl;
  wire swap_1_nor_1_nl;
  wire swap_1_swap_1_and_9_nl;
  wire while_if_while_if_nor_67_nl;
  wire low_or_nl;
  wire[32:0] while_acc_3_nl;
  wire[33:0] nl_while_acc_3_nl;
  wire[33:0] acc_nl;
  wire[34:0] nl_acc_nl;
  wire[1:0] while_and_250_nl;
  wire[1:0] while_mux1h_3_nl;
  wire while_nor_3_nl;
  wire[29:0] while_mux1h_4_nl;
  wire while_or_196_nl;
  wire[31:0] while_while_while_nand_1_nl;
  wire[31:0] while_mux_1_nl;
  wire while_nor_5_nl;
  wire[33:0] acc_1_nl;
  wire[34:0] nl_acc_1_nl;
  wire[31:0] partition_while_while_mux_5_nl;
  wire[5:0] partition_pivot_mux1h_71_nl;
  wire or_798_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_arr_rsci_ldout;
  assign nl_arr_rsci_ldout = ((z_out_1[32]) & (fsm_output[6])) | (while_acc_3_cse_32
      & (fsm_output[8]));
  wire[31:0] partition_pivot_partition_pivot_mux1h_63_nl;
  wire partition_pivot_or_126_nl;
  wire partition_pivot_or_127_nl;
  wire partition_pivot_or_128_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_62_nl;
  wire partition_pivot_or_124_nl;
  wire partition_pivot_or_125_nl;
  wire partition_pivot_or_129_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_61_nl;
  wire partition_pivot_or_122_nl;
  wire partition_pivot_or_123_nl;
  wire partition_pivot_or_130_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_60_nl;
  wire partition_pivot_or_120_nl;
  wire partition_pivot_or_121_nl;
  wire partition_pivot_or_131_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_59_nl;
  wire partition_pivot_or_118_nl;
  wire partition_pivot_or_119_nl;
  wire partition_pivot_or_132_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_58_nl;
  wire partition_pivot_or_116_nl;
  wire partition_pivot_or_117_nl;
  wire partition_pivot_or_133_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_57_nl;
  wire partition_pivot_or_114_nl;
  wire partition_pivot_or_115_nl;
  wire partition_pivot_or_134_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_56_nl;
  wire partition_pivot_or_112_nl;
  wire partition_pivot_or_113_nl;
  wire partition_pivot_or_135_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_55_nl;
  wire partition_pivot_or_110_nl;
  wire partition_pivot_or_111_nl;
  wire partition_pivot_or_136_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_54_nl;
  wire partition_pivot_or_108_nl;
  wire partition_pivot_or_109_nl;
  wire partition_pivot_or_137_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_53_nl;
  wire partition_pivot_or_106_nl;
  wire partition_pivot_or_107_nl;
  wire partition_pivot_or_138_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_52_nl;
  wire partition_pivot_or_104_nl;
  wire partition_pivot_or_105_nl;
  wire partition_pivot_or_139_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_51_nl;
  wire partition_pivot_or_102_nl;
  wire partition_pivot_or_103_nl;
  wire partition_pivot_or_140_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_50_nl;
  wire partition_pivot_or_100_nl;
  wire partition_pivot_or_101_nl;
  wire partition_pivot_or_141_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_49_nl;
  wire partition_pivot_or_98_nl;
  wire partition_pivot_or_99_nl;
  wire partition_pivot_or_142_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_48_nl;
  wire partition_pivot_or_96_nl;
  wire partition_pivot_or_97_nl;
  wire partition_pivot_or_143_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_47_nl;
  wire partition_pivot_or_94_nl;
  wire partition_pivot_or_95_nl;
  wire partition_pivot_or_144_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_46_nl;
  wire partition_pivot_or_92_nl;
  wire partition_pivot_or_93_nl;
  wire partition_pivot_or_145_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_45_nl;
  wire partition_pivot_or_90_nl;
  wire partition_pivot_or_91_nl;
  wire partition_pivot_or_146_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_44_nl;
  wire partition_pivot_or_88_nl;
  wire partition_pivot_or_89_nl;
  wire partition_pivot_or_147_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_43_nl;
  wire partition_pivot_or_86_nl;
  wire partition_pivot_or_87_nl;
  wire partition_pivot_or_148_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_42_nl;
  wire partition_pivot_or_84_nl;
  wire partition_pivot_or_85_nl;
  wire partition_pivot_or_149_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_41_nl;
  wire partition_pivot_or_82_nl;
  wire partition_pivot_or_83_nl;
  wire partition_pivot_or_150_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_40_nl;
  wire partition_pivot_or_80_nl;
  wire partition_pivot_or_81_nl;
  wire partition_pivot_or_151_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_39_nl;
  wire partition_pivot_or_78_nl;
  wire partition_pivot_or_79_nl;
  wire partition_pivot_or_152_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_38_nl;
  wire partition_pivot_or_76_nl;
  wire partition_pivot_or_77_nl;
  wire partition_pivot_or_153_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_37_nl;
  wire partition_pivot_or_74_nl;
  wire partition_pivot_or_75_nl;
  wire partition_pivot_or_154_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_36_nl;
  wire partition_pivot_or_72_nl;
  wire partition_pivot_or_73_nl;
  wire partition_pivot_or_155_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_35_nl;
  wire partition_pivot_or_70_nl;
  wire partition_pivot_or_71_nl;
  wire partition_pivot_or_156_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_34_nl;
  wire partition_pivot_or_68_nl;
  wire partition_pivot_or_69_nl;
  wire partition_pivot_or_157_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_33_nl;
  wire partition_pivot_or_66_nl;
  wire partition_pivot_or_67_nl;
  wire partition_pivot_or_158_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_32_nl;
  wire partition_pivot_or_64_nl;
  wire partition_pivot_or_65_nl;
  wire partition_pivot_or_159_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_31_nl;
  wire partition_pivot_or_62_nl;
  wire partition_pivot_or_63_nl;
  wire partition_pivot_or_160_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_30_nl;
  wire partition_pivot_or_60_nl;
  wire partition_pivot_or_61_nl;
  wire partition_pivot_or_161_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_29_nl;
  wire partition_pivot_or_58_nl;
  wire partition_pivot_or_59_nl;
  wire partition_pivot_or_162_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_28_nl;
  wire partition_pivot_or_56_nl;
  wire partition_pivot_or_57_nl;
  wire partition_pivot_or_163_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_27_nl;
  wire partition_pivot_or_54_nl;
  wire partition_pivot_or_55_nl;
  wire partition_pivot_or_164_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_26_nl;
  wire partition_pivot_or_52_nl;
  wire partition_pivot_or_53_nl;
  wire partition_pivot_or_165_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_25_nl;
  wire partition_pivot_or_50_nl;
  wire partition_pivot_or_51_nl;
  wire partition_pivot_or_166_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_24_nl;
  wire partition_pivot_or_48_nl;
  wire partition_pivot_or_49_nl;
  wire partition_pivot_or_167_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_23_nl;
  wire partition_pivot_or_46_nl;
  wire partition_pivot_or_47_nl;
  wire partition_pivot_or_168_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_22_nl;
  wire partition_pivot_or_44_nl;
  wire partition_pivot_or_45_nl;
  wire partition_pivot_or_169_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_21_nl;
  wire partition_pivot_or_42_nl;
  wire partition_pivot_or_43_nl;
  wire partition_pivot_or_170_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_20_nl;
  wire partition_pivot_or_40_nl;
  wire partition_pivot_or_41_nl;
  wire partition_pivot_or_171_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_19_nl;
  wire partition_pivot_or_38_nl;
  wire partition_pivot_or_39_nl;
  wire partition_pivot_or_172_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_18_nl;
  wire partition_pivot_or_36_nl;
  wire partition_pivot_or_37_nl;
  wire partition_pivot_or_173_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_17_nl;
  wire partition_pivot_or_34_nl;
  wire partition_pivot_or_35_nl;
  wire partition_pivot_or_174_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_16_nl;
  wire partition_pivot_or_32_nl;
  wire partition_pivot_or_33_nl;
  wire partition_pivot_or_175_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_15_nl;
  wire partition_pivot_or_30_nl;
  wire partition_pivot_or_31_nl;
  wire partition_pivot_or_176_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_14_nl;
  wire partition_pivot_or_28_nl;
  wire partition_pivot_or_29_nl;
  wire partition_pivot_or_177_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_13_nl;
  wire partition_pivot_or_26_nl;
  wire partition_pivot_or_27_nl;
  wire partition_pivot_or_178_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_12_nl;
  wire partition_pivot_or_24_nl;
  wire partition_pivot_or_25_nl;
  wire partition_pivot_or_179_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_11_nl;
  wire partition_pivot_or_22_nl;
  wire partition_pivot_or_23_nl;
  wire partition_pivot_or_180_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_10_nl;
  wire partition_pivot_or_20_nl;
  wire partition_pivot_or_21_nl;
  wire partition_pivot_or_181_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_9_nl;
  wire partition_pivot_or_18_nl;
  wire partition_pivot_or_19_nl;
  wire partition_pivot_or_182_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_8_nl;
  wire partition_pivot_or_16_nl;
  wire partition_pivot_or_17_nl;
  wire partition_pivot_or_183_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_7_nl;
  wire partition_pivot_or_14_nl;
  wire partition_pivot_or_15_nl;
  wire partition_pivot_or_184_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_6_nl;
  wire partition_pivot_or_12_nl;
  wire partition_pivot_or_13_nl;
  wire partition_pivot_or_185_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_5_nl;
  wire partition_pivot_or_10_nl;
  wire partition_pivot_or_11_nl;
  wire partition_pivot_or_186_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_4_nl;
  wire partition_pivot_or_8_nl;
  wire partition_pivot_or_9_nl;
  wire partition_pivot_or_187_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_3_nl;
  wire partition_pivot_or_6_nl;
  wire partition_pivot_or_7_nl;
  wire partition_pivot_or_188_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_2_nl;
  wire partition_pivot_or_4_nl;
  wire partition_pivot_or_5_nl;
  wire partition_pivot_or_189_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_1_nl;
  wire partition_pivot_or_2_nl;
  wire partition_pivot_or_3_nl;
  wire partition_pivot_or_190_nl;
  wire[31:0] partition_pivot_partition_pivot_mux1h_nl;
  wire partition_pivot_or_191_nl;
  wire partition_pivot_or_nl;
  wire partition_pivot_or_1_nl;
  wire [2047:0] nl_arr_rsci_dout;
  assign partition_pivot_or_126_nl = (~(swap_equal_tmp_176 | swap_equal_tmp_128 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_63 | swap_1_equal_tmp_127)) & (fsm_output[8]));
  assign partition_pivot_or_127_nl = (swap_equal_tmp_176 & (~ swap_equal_tmp_128)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_63 & (~ swap_1_equal_tmp_127) &
      (fsm_output[8]));
  assign partition_pivot_or_128_nl = (swap_equal_tmp_128 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_127 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_63_nl = MUX1HOT_v_32_3_2((arr_rsci_din[2047:2016]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_126_nl , partition_pivot_or_127_nl
      , partition_pivot_or_128_nl});
  assign partition_pivot_or_124_nl = (~(swap_equal_tmp_177 | swap_equal_tmp_129 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_62 | swap_1_equal_tmp_126)) & (fsm_output[8]));
  assign partition_pivot_or_125_nl = (swap_equal_tmp_177 & (~ swap_equal_tmp_129)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_62 & (~ swap_1_equal_tmp_126) &
      (fsm_output[8]));
  assign partition_pivot_or_129_nl = (swap_equal_tmp_129 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_126 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_62_nl = MUX1HOT_v_32_3_2((arr_rsci_din[2015:1984]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_124_nl , partition_pivot_or_125_nl
      , partition_pivot_or_129_nl});
  assign partition_pivot_or_122_nl = (~(swap_equal_tmp_180 | swap_equal_tmp_130 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_61 | swap_1_equal_tmp_125)) & (fsm_output[8]));
  assign partition_pivot_or_123_nl = (swap_equal_tmp_180 & (~ swap_equal_tmp_130)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_61 & (~ swap_1_equal_tmp_125) &
      (fsm_output[8]));
  assign partition_pivot_or_130_nl = (swap_equal_tmp_130 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_125 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_61_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1983:1952]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_122_nl , partition_pivot_or_123_nl
      , partition_pivot_or_130_nl});
  assign partition_pivot_or_120_nl = (~(swap_equal_tmp_183 | swap_equal_tmp_131 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_60 | swap_1_equal_tmp_124)) & (fsm_output[8]));
  assign partition_pivot_or_121_nl = (swap_equal_tmp_183 & (~ swap_equal_tmp_131)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_60 & (~ swap_1_equal_tmp_124) &
      (fsm_output[8]));
  assign partition_pivot_or_131_nl = (swap_equal_tmp_131 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_124 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_60_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1951:1920]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_120_nl , partition_pivot_or_121_nl
      , partition_pivot_or_131_nl});
  assign partition_pivot_or_118_nl = (~(swap_equal_tmp_186 | swap_equal_tmp_132 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_59 | swap_1_equal_tmp_123)) & (fsm_output[8]));
  assign partition_pivot_or_119_nl = (swap_equal_tmp_186 & (~ swap_equal_tmp_132)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_59 & (~ swap_1_equal_tmp_123) &
      (fsm_output[8]));
  assign partition_pivot_or_132_nl = (swap_equal_tmp_132 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_123 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_59_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1919:1888]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_118_nl , partition_pivot_or_119_nl
      , partition_pivot_or_132_nl});
  assign partition_pivot_or_116_nl = (~(swap_equal_tmp_189 | swap_equal_tmp_133 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_58 | swap_1_equal_tmp_122)) & (fsm_output[8]));
  assign partition_pivot_or_117_nl = (swap_equal_tmp_189 & (~ swap_equal_tmp_133)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_58 & (~ swap_1_equal_tmp_122) &
      (fsm_output[8]));
  assign partition_pivot_or_133_nl = (swap_equal_tmp_133 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_122 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_58_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1887:1856]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_116_nl , partition_pivot_or_117_nl
      , partition_pivot_or_133_nl});
  assign partition_pivot_or_114_nl = (~(swap_equal_tmp_192 | swap_equal_tmp_134 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_57 | swap_1_equal_tmp_121)) & (fsm_output[8]));
  assign partition_pivot_or_115_nl = (swap_equal_tmp_192 & (~ swap_equal_tmp_134)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_57 & (~ swap_1_equal_tmp_121) &
      (fsm_output[8]));
  assign partition_pivot_or_134_nl = (swap_equal_tmp_134 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_121 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_57_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1855:1824]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_114_nl , partition_pivot_or_115_nl
      , partition_pivot_or_134_nl});
  assign partition_pivot_or_112_nl = (~(swap_equal_tmp_195 | swap_equal_tmp_135 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_56 | swap_1_equal_tmp_120)) & (fsm_output[8]));
  assign partition_pivot_or_113_nl = (swap_equal_tmp_195 & (~ swap_equal_tmp_135)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_56 & (~ swap_1_equal_tmp_120) &
      (fsm_output[8]));
  assign partition_pivot_or_135_nl = (swap_equal_tmp_135 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_120 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_56_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1823:1792]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_112_nl , partition_pivot_or_113_nl
      , partition_pivot_or_135_nl});
  assign partition_pivot_or_110_nl = (~(swap_equal_tmp_197 | swap_equal_tmp_137 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_55 | swap_1_equal_tmp_119)) & (fsm_output[8]));
  assign partition_pivot_or_111_nl = (swap_equal_tmp_197 & (~ swap_equal_tmp_137)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_55 & (~ swap_1_equal_tmp_119) &
      (fsm_output[8]));
  assign partition_pivot_or_136_nl = (swap_equal_tmp_137 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_119 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_55_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1791:1760]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_110_nl , partition_pivot_or_111_nl
      , partition_pivot_or_136_nl});
  assign partition_pivot_or_108_nl = (~(swap_equal_tmp_200 | swap_equal_tmp_138 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_54 | swap_1_equal_tmp_118)) & (fsm_output[8]));
  assign partition_pivot_or_109_nl = (swap_equal_tmp_200 & (~ swap_equal_tmp_138)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_54 & (~ swap_1_equal_tmp_118) &
      (fsm_output[8]));
  assign partition_pivot_or_137_nl = (swap_equal_tmp_138 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_118 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_54_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1759:1728]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_108_nl , partition_pivot_or_109_nl
      , partition_pivot_or_137_nl});
  assign partition_pivot_or_106_nl = (~(swap_equal_tmp_202 | swap_equal_tmp_140 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_53 | swap_1_equal_tmp_117)) & (fsm_output[8]));
  assign partition_pivot_or_107_nl = (swap_equal_tmp_202 & (~ swap_equal_tmp_140)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_53 & (~ swap_1_equal_tmp_117) &
      (fsm_output[8]));
  assign partition_pivot_or_138_nl = (swap_equal_tmp_140 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_117 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_53_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1727:1696]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_106_nl , partition_pivot_or_107_nl
      , partition_pivot_or_138_nl});
  assign partition_pivot_or_104_nl = (~(swap_equal_tmp_204 | swap_equal_tmp_142 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_52 | swap_1_equal_tmp_116)) & (fsm_output[8]));
  assign partition_pivot_or_105_nl = (swap_equal_tmp_204 & (~ swap_equal_tmp_142)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_52 & (~ swap_1_equal_tmp_116) &
      (fsm_output[8]));
  assign partition_pivot_or_139_nl = (swap_equal_tmp_142 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_116 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_52_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1695:1664]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_104_nl , partition_pivot_or_105_nl
      , partition_pivot_or_139_nl});
  assign partition_pivot_or_102_nl = (~(swap_equal_tmp_206 | swap_equal_tmp_144 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_51 | swap_1_equal_tmp_115)) & (fsm_output[8]));
  assign partition_pivot_or_103_nl = (swap_equal_tmp_206 & (~ swap_equal_tmp_144)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_51 & (~ swap_1_equal_tmp_115) &
      (fsm_output[8]));
  assign partition_pivot_or_140_nl = (swap_equal_tmp_144 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_115 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_51_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1663:1632]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_102_nl , partition_pivot_or_103_nl
      , partition_pivot_or_140_nl});
  assign partition_pivot_or_100_nl = (~(swap_equal_tmp_208 | swap_equal_tmp_146 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_50 | swap_1_equal_tmp_114)) & (fsm_output[8]));
  assign partition_pivot_or_101_nl = (swap_equal_tmp_208 & (~ swap_equal_tmp_146)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_50 & (~ swap_1_equal_tmp_114) &
      (fsm_output[8]));
  assign partition_pivot_or_141_nl = (swap_equal_tmp_146 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_114 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_50_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1631:1600]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_100_nl , partition_pivot_or_101_nl
      , partition_pivot_or_141_nl});
  assign partition_pivot_or_98_nl = (~(swap_equal_tmp_210 | swap_equal_tmp_148 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_49 | swap_1_equal_tmp_113)) & (fsm_output[8]));
  assign partition_pivot_or_99_nl = (swap_equal_tmp_210 & (~ swap_equal_tmp_148)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_49 & (~ swap_1_equal_tmp_113) &
      (fsm_output[8]));
  assign partition_pivot_or_142_nl = (swap_equal_tmp_148 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_113 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_49_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1599:1568]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_98_nl , partition_pivot_or_99_nl
      , partition_pivot_or_142_nl});
  assign partition_pivot_or_96_nl = (~(swap_equal_tmp_212 | swap_equal_tmp_213 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_48 | swap_1_equal_tmp_297)) & (fsm_output[8]));
  assign partition_pivot_or_97_nl = (swap_equal_tmp_212 & (~ swap_equal_tmp_213)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_48 & (~ swap_1_equal_tmp_297) &
      (fsm_output[8]));
  assign partition_pivot_or_143_nl = (swap_equal_tmp_213 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_297 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_48_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1567:1536]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_96_nl , partition_pivot_or_97_nl
      , partition_pivot_or_143_nl});
  assign partition_pivot_or_94_nl = (~(swap_equal_tmp_215 | swap_equal_tmp_151 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_47 | swap_1_equal_tmp_111)) & (fsm_output[8]));
  assign partition_pivot_or_95_nl = (swap_equal_tmp_215 & (~ swap_equal_tmp_151)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_47 & (~ swap_1_equal_tmp_111) &
      (fsm_output[8]));
  assign partition_pivot_or_144_nl = (swap_equal_tmp_151 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_111 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_47_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1535:1504]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_94_nl , partition_pivot_or_95_nl
      , partition_pivot_or_144_nl});
  assign partition_pivot_or_92_nl = (~(swap_equal_tmp_218 | swap_equal_tmp_152 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_46 | swap_1_equal_tmp_110)) & (fsm_output[8]));
  assign partition_pivot_or_93_nl = (swap_equal_tmp_218 & (~ swap_equal_tmp_152)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_46 & (~ swap_1_equal_tmp_110) &
      (fsm_output[8]));
  assign partition_pivot_or_145_nl = (swap_equal_tmp_152 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_110 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_46_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1503:1472]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_92_nl , partition_pivot_or_93_nl
      , partition_pivot_or_145_nl});
  assign partition_pivot_or_90_nl = (~(swap_equal_tmp_221 | swap_equal_tmp_153 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_45 | swap_1_equal_tmp_109)) & (fsm_output[8]));
  assign partition_pivot_or_91_nl = (swap_equal_tmp_221 & (~ swap_equal_tmp_153)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_45 & (~ swap_1_equal_tmp_109) &
      (fsm_output[8]));
  assign partition_pivot_or_146_nl = (swap_equal_tmp_153 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_109 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_45_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1471:1440]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_90_nl , partition_pivot_or_91_nl
      , partition_pivot_or_146_nl});
  assign partition_pivot_or_88_nl = (~(swap_equal_tmp_224 | swap_equal_tmp_154 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_44 | swap_1_equal_tmp_108)) & (fsm_output[8]));
  assign partition_pivot_or_89_nl = (swap_equal_tmp_224 & (~ swap_equal_tmp_154)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_44 & (~ swap_1_equal_tmp_108) &
      (fsm_output[8]));
  assign partition_pivot_or_147_nl = (swap_equal_tmp_154 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_108 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_44_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1439:1408]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_88_nl , partition_pivot_or_89_nl
      , partition_pivot_or_147_nl});
  assign partition_pivot_or_86_nl = (~(swap_equal_tmp_226 | swap_equal_tmp_156 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_43 | swap_1_equal_tmp_107)) & (fsm_output[8]));
  assign partition_pivot_or_87_nl = (swap_equal_tmp_226 & (~ swap_equal_tmp_156)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_43 & (~ swap_1_equal_tmp_107) &
      (fsm_output[8]));
  assign partition_pivot_or_148_nl = (swap_equal_tmp_156 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_107 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_43_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1407:1376]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_86_nl , partition_pivot_or_87_nl
      , partition_pivot_or_148_nl});
  assign partition_pivot_or_84_nl = (~(swap_equal_tmp_229 | swap_equal_tmp_157 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_42 | swap_1_equal_tmp_106)) & (fsm_output[8]));
  assign partition_pivot_or_85_nl = (swap_equal_tmp_229 & (~ swap_equal_tmp_157)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_42 & (~ swap_1_equal_tmp_106) &
      (fsm_output[8]));
  assign partition_pivot_or_149_nl = (swap_equal_tmp_157 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_106 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_42_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1375:1344]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_84_nl , partition_pivot_or_85_nl
      , partition_pivot_or_149_nl});
  assign partition_pivot_or_82_nl = (~(swap_equal_tmp_231 | swap_equal_tmp_159 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_41 | swap_1_equal_tmp_105)) & (fsm_output[8]));
  assign partition_pivot_or_83_nl = (swap_equal_tmp_231 & (~ swap_equal_tmp_159)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_41 & (~ swap_1_equal_tmp_105) &
      (fsm_output[8]));
  assign partition_pivot_or_150_nl = (swap_equal_tmp_159 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_105 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_41_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1343:1312]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_82_nl , partition_pivot_or_83_nl
      , partition_pivot_or_150_nl});
  assign partition_pivot_or_80_nl = (~(swap_equal_tmp_233 | swap_equal_tmp_234 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_40 | swap_1_equal_tmp_303)) & (fsm_output[8]));
  assign partition_pivot_or_81_nl = (swap_equal_tmp_233 & (~ swap_equal_tmp_234)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_40 & (~ swap_1_equal_tmp_303) &
      (fsm_output[8]));
  assign partition_pivot_or_151_nl = (swap_equal_tmp_234 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_303 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_40_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1311:1280]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_80_nl , partition_pivot_or_81_nl
      , partition_pivot_or_151_nl});
  assign partition_pivot_or_78_nl = (~(swap_equal_tmp_236 | swap_equal_tmp_162 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_39 | swap_1_equal_tmp_103)) & (fsm_output[8]));
  assign partition_pivot_or_79_nl = (swap_equal_tmp_236 & (~ swap_equal_tmp_162)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_39 & (~ swap_1_equal_tmp_103) &
      (fsm_output[8]));
  assign partition_pivot_or_152_nl = (swap_equal_tmp_162 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_103 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_39_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1279:1248]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_78_nl , partition_pivot_or_79_nl
      , partition_pivot_or_152_nl});
  assign partition_pivot_or_76_nl = (~(swap_equal_tmp_238 | swap_equal_tmp_164 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_38 | swap_1_equal_tmp_102)) & (fsm_output[8]));
  assign partition_pivot_or_77_nl = (swap_equal_tmp_238 & (~ swap_equal_tmp_164)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_38 & (~ swap_1_equal_tmp_102) &
      (fsm_output[8]));
  assign partition_pivot_or_153_nl = (swap_equal_tmp_164 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_102 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_38_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1247:1216]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_76_nl , partition_pivot_or_77_nl
      , partition_pivot_or_153_nl});
  assign partition_pivot_or_74_nl = (~(swap_equal_tmp_240 | swap_equal_tmp_166 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_37 | swap_1_equal_tmp_101)) & (fsm_output[8]));
  assign partition_pivot_or_75_nl = (swap_equal_tmp_240 & (~ swap_equal_tmp_166)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_37 & (~ swap_1_equal_tmp_101) &
      (fsm_output[8]));
  assign partition_pivot_or_154_nl = (swap_equal_tmp_166 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_101 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_37_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1215:1184]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_74_nl , partition_pivot_or_75_nl
      , partition_pivot_or_154_nl});
  assign partition_pivot_or_72_nl = (~(swap_equal_tmp_242 | swap_equal_tmp_168 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_36 | swap_1_equal_tmp_100)) & (fsm_output[8]));
  assign partition_pivot_or_73_nl = (swap_equal_tmp_242 & (~ swap_equal_tmp_168)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_36 & (~ swap_1_equal_tmp_100) &
      (fsm_output[8]));
  assign partition_pivot_or_155_nl = (swap_equal_tmp_168 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_100 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_36_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1183:1152]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_72_nl , partition_pivot_or_73_nl
      , partition_pivot_or_155_nl});
  assign partition_pivot_or_70_nl = (~(swap_equal_tmp_244 | swap_equal_tmp_170 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_35 | swap_1_equal_tmp_99)) & (fsm_output[8]));
  assign partition_pivot_or_71_nl = (swap_equal_tmp_244 & (~ swap_equal_tmp_170)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_35 & (~ swap_1_equal_tmp_99) & (fsm_output[8]));
  assign partition_pivot_or_156_nl = (swap_equal_tmp_170 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_99 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_35_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1151:1120]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_70_nl , partition_pivot_or_71_nl
      , partition_pivot_or_156_nl});
  assign partition_pivot_or_68_nl = (~(swap_equal_tmp_246 | swap_equal_tmp_247 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_34 | swap_1_equal_tmp_304)) & (fsm_output[8]));
  assign partition_pivot_or_69_nl = (swap_equal_tmp_246 & (~ swap_equal_tmp_247)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_34 & (~ swap_1_equal_tmp_304) &
      (fsm_output[8]));
  assign partition_pivot_or_157_nl = (swap_equal_tmp_247 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_304 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_34_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1119:1088]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_68_nl , partition_pivot_or_69_nl
      , partition_pivot_or_157_nl});
  assign partition_pivot_or_66_nl = (~(swap_equal_tmp_249 | swap_equal_tmp_173 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_33 | swap_1_equal_tmp_97)) & (fsm_output[8]));
  assign partition_pivot_or_67_nl = (swap_equal_tmp_249 & (~ swap_equal_tmp_173)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_33 & (~ swap_1_equal_tmp_97) & (fsm_output[8]));
  assign partition_pivot_or_158_nl = (swap_equal_tmp_173 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_97 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_33_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1087:1056]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_66_nl , partition_pivot_or_67_nl
      , partition_pivot_or_158_nl});
  assign partition_pivot_or_64_nl = (~(swap_equal_tmp_251 | swap_equal_tmp_252 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_305 | swap_1_equal_tmp_306)) & (fsm_output[8]));
  assign partition_pivot_or_65_nl = (swap_equal_tmp_251 & (~ swap_equal_tmp_252)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_305 & (~ swap_1_equal_tmp_306) &
      (fsm_output[8]));
  assign partition_pivot_or_159_nl = (swap_equal_tmp_252 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_306 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_32_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1055:1024]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_64_nl , partition_pivot_or_65_nl
      , partition_pivot_or_159_nl});
  assign partition_pivot_or_62_nl = (~(swap_equal_tmp_253 | swap_equal_tmp_175 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_31 | swap_1_equal_tmp_95)) & (fsm_output[8]));
  assign partition_pivot_or_63_nl = (swap_equal_tmp_253 & (~ swap_equal_tmp_175)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_31 & (~ swap_1_equal_tmp_95) & (fsm_output[8]));
  assign partition_pivot_or_160_nl = (swap_equal_tmp_175 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_95 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_31_nl = MUX1HOT_v_32_3_2((arr_rsci_din[1023:992]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_62_nl , partition_pivot_or_63_nl
      , partition_pivot_or_160_nl});
  assign partition_pivot_or_60_nl = (~(swap_equal_tmp_250 | swap_equal_tmp_174 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_30 | swap_1_equal_tmp_94)) & (fsm_output[8]));
  assign partition_pivot_or_61_nl = (swap_equal_tmp_250 & (~ swap_equal_tmp_174)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_30 & (~ swap_1_equal_tmp_94) & (fsm_output[8]));
  assign partition_pivot_or_161_nl = (swap_equal_tmp_174 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_94 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_30_nl = MUX1HOT_v_32_3_2((arr_rsci_din[991:960]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_60_nl , partition_pivot_or_61_nl
      , partition_pivot_or_161_nl});
  assign partition_pivot_or_58_nl = (~(swap_equal_tmp_248 | swap_equal_tmp_172 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_29 | swap_1_equal_tmp_93)) & (fsm_output[8]));
  assign partition_pivot_or_59_nl = (swap_equal_tmp_248 & (~ swap_equal_tmp_172)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_29 & (~ swap_1_equal_tmp_93) & (fsm_output[8]));
  assign partition_pivot_or_162_nl = (swap_equal_tmp_172 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_93 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_29_nl = MUX1HOT_v_32_3_2((arr_rsci_din[959:928]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_58_nl , partition_pivot_or_59_nl
      , partition_pivot_or_162_nl});
  assign partition_pivot_or_56_nl = (~(swap_equal_tmp_245 | swap_equal_tmp_171 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_28 | swap_1_equal_tmp_92)) & (fsm_output[8]));
  assign partition_pivot_or_57_nl = (swap_equal_tmp_245 & (~ swap_equal_tmp_171)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_28 & (~ swap_1_equal_tmp_92) & (fsm_output[8]));
  assign partition_pivot_or_163_nl = (swap_equal_tmp_171 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_92 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_28_nl = MUX1HOT_v_32_3_2((arr_rsci_din[927:896]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_56_nl , partition_pivot_or_57_nl
      , partition_pivot_or_163_nl});
  assign partition_pivot_or_54_nl = (~(swap_equal_tmp_243 | swap_equal_tmp_169 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_27 | swap_1_equal_tmp_91)) & (fsm_output[8]));
  assign partition_pivot_or_55_nl = (swap_equal_tmp_243 & (~ swap_equal_tmp_169)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_27 & (~ swap_1_equal_tmp_91) & (fsm_output[8]));
  assign partition_pivot_or_164_nl = (swap_equal_tmp_169 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_91 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_27_nl = MUX1HOT_v_32_3_2((arr_rsci_din[895:864]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_54_nl , partition_pivot_or_55_nl
      , partition_pivot_or_164_nl});
  assign partition_pivot_or_52_nl = (~(swap_equal_tmp_241 | swap_equal_tmp_167 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_26 | swap_1_equal_tmp_90)) & (fsm_output[8]));
  assign partition_pivot_or_53_nl = (swap_equal_tmp_241 & (~ swap_equal_tmp_167)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_26 & (~ swap_1_equal_tmp_90) & (fsm_output[8]));
  assign partition_pivot_or_165_nl = (swap_equal_tmp_167 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_90 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_26_nl = MUX1HOT_v_32_3_2((arr_rsci_din[863:832]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_52_nl , partition_pivot_or_53_nl
      , partition_pivot_or_165_nl});
  assign partition_pivot_or_50_nl = (~(swap_equal_tmp_239 | swap_equal_tmp_165 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_25 | swap_1_equal_tmp_89)) & (fsm_output[8]));
  assign partition_pivot_or_51_nl = (swap_equal_tmp_239 & (~ swap_equal_tmp_165)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_25 & (~ swap_1_equal_tmp_89) & (fsm_output[8]));
  assign partition_pivot_or_166_nl = (swap_equal_tmp_165 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_89 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_25_nl = MUX1HOT_v_32_3_2((arr_rsci_din[831:800]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_50_nl , partition_pivot_or_51_nl
      , partition_pivot_or_166_nl});
  assign partition_pivot_or_48_nl = (~(swap_equal_tmp_237 | swap_equal_tmp_163 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_24 | swap_1_equal_tmp_88)) & (fsm_output[8]));
  assign partition_pivot_or_49_nl = (swap_equal_tmp_237 & (~ swap_equal_tmp_163)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_24 & (~ swap_1_equal_tmp_88) & (fsm_output[8]));
  assign partition_pivot_or_167_nl = (swap_equal_tmp_163 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_88 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_24_nl = MUX1HOT_v_32_3_2((arr_rsci_din[799:768]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_48_nl , partition_pivot_or_49_nl
      , partition_pivot_or_167_nl});
  assign partition_pivot_or_46_nl = (~(swap_equal_tmp_235 | swap_equal_tmp_161 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_23 | swap_1_equal_tmp_87)) & (fsm_output[8]));
  assign partition_pivot_or_47_nl = (swap_equal_tmp_235 & (~ swap_equal_tmp_161)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_23 & (~ swap_1_equal_tmp_87) & (fsm_output[8]));
  assign partition_pivot_or_168_nl = (swap_equal_tmp_161 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_87 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_23_nl = MUX1HOT_v_32_3_2((arr_rsci_din[767:736]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_46_nl , partition_pivot_or_47_nl
      , partition_pivot_or_168_nl});
  assign partition_pivot_or_44_nl = (~(swap_equal_tmp_232 | swap_equal_tmp_160 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_22 | swap_1_equal_tmp_86)) & (fsm_output[8]));
  assign partition_pivot_or_45_nl = (swap_equal_tmp_232 & (~ swap_equal_tmp_160)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_22 & (~ swap_1_equal_tmp_86) & (fsm_output[8]));
  assign partition_pivot_or_169_nl = (swap_equal_tmp_160 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_86 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_22_nl = MUX1HOT_v_32_3_2((arr_rsci_din[735:704]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_44_nl , partition_pivot_or_45_nl
      , partition_pivot_or_169_nl});
  assign partition_pivot_or_42_nl = (~(swap_equal_tmp_230 | swap_equal_tmp_158 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_21 | swap_1_equal_tmp_85)) & (fsm_output[8]));
  assign partition_pivot_or_43_nl = (swap_equal_tmp_230 & (~ swap_equal_tmp_158)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_21 & (~ swap_1_equal_tmp_85) & (fsm_output[8]));
  assign partition_pivot_or_170_nl = (swap_equal_tmp_158 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_85 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_21_nl = MUX1HOT_v_32_3_2((arr_rsci_din[703:672]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_42_nl , partition_pivot_or_43_nl
      , partition_pivot_or_170_nl});
  assign partition_pivot_or_40_nl = (~(swap_equal_tmp_227 | swap_equal_tmp_228 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_20 | swap_1_equal_tmp_302)) & (fsm_output[8]));
  assign partition_pivot_or_41_nl = (swap_equal_tmp_227 & (~ swap_equal_tmp_228)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_20 & (~ swap_1_equal_tmp_302) &
      (fsm_output[8]));
  assign partition_pivot_or_171_nl = (swap_equal_tmp_228 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_302 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_20_nl = MUX1HOT_v_32_3_2((arr_rsci_din[671:640]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_40_nl , partition_pivot_or_41_nl
      , partition_pivot_or_171_nl});
  assign partition_pivot_or_38_nl = (~(swap_equal_tmp_225 | swap_equal_tmp_155 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_19 | swap_1_equal_tmp_83)) & (fsm_output[8]));
  assign partition_pivot_or_39_nl = (swap_equal_tmp_225 & (~ swap_equal_tmp_155)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_19 & (~ swap_1_equal_tmp_83) & (fsm_output[8]));
  assign partition_pivot_or_172_nl = (swap_equal_tmp_155 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_83 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_19_nl = MUX1HOT_v_32_3_2((arr_rsci_din[639:608]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_38_nl , partition_pivot_or_39_nl
      , partition_pivot_or_172_nl});
  assign partition_pivot_or_36_nl = (~(swap_equal_tmp_222 | swap_equal_tmp_223 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_18 | swap_1_equal_tmp_301)) & (fsm_output[8]));
  assign partition_pivot_or_37_nl = (swap_equal_tmp_222 & (~ swap_equal_tmp_223)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_18 & (~ swap_1_equal_tmp_301) &
      (fsm_output[8]));
  assign partition_pivot_or_173_nl = (swap_equal_tmp_223 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_301 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_18_nl = MUX1HOT_v_32_3_2((arr_rsci_din[607:576]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_36_nl , partition_pivot_or_37_nl
      , partition_pivot_or_173_nl});
  assign partition_pivot_or_34_nl = (~(swap_equal_tmp_219 | swap_equal_tmp_220 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_17 | swap_1_equal_tmp_300)) & (fsm_output[8]));
  assign partition_pivot_or_35_nl = (swap_equal_tmp_219 & (~ swap_equal_tmp_220)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_17 & (~ swap_1_equal_tmp_300) &
      (fsm_output[8]));
  assign partition_pivot_or_174_nl = (swap_equal_tmp_220 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_300 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_17_nl = MUX1HOT_v_32_3_2((arr_rsci_din[575:544]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_34_nl , partition_pivot_or_35_nl
      , partition_pivot_or_174_nl});
  assign partition_pivot_or_32_nl = (~(swap_equal_tmp_216 | swap_equal_tmp_217 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_298 | swap_1_equal_tmp_299)) & (fsm_output[8]));
  assign partition_pivot_or_33_nl = (swap_equal_tmp_216 & (~ swap_equal_tmp_217)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_298 & (~ swap_1_equal_tmp_299) &
      (fsm_output[8]));
  assign partition_pivot_or_175_nl = (swap_equal_tmp_217 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_299 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_16_nl = MUX1HOT_v_32_3_2((arr_rsci_din[543:512]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_32_nl , partition_pivot_or_33_nl
      , partition_pivot_or_175_nl});
  assign partition_pivot_or_30_nl = (~(swap_equal_tmp_214 | swap_equal_tmp_150 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_15 | swap_1_equal_tmp_79)) & (fsm_output[8]));
  assign partition_pivot_or_31_nl = (swap_equal_tmp_214 & (~ swap_equal_tmp_150)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_15 & (~ swap_1_equal_tmp_79) & (fsm_output[8]));
  assign partition_pivot_or_176_nl = (swap_equal_tmp_150 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_79 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_15_nl = MUX1HOT_v_32_3_2((arr_rsci_din[511:480]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_30_nl , partition_pivot_or_31_nl
      , partition_pivot_or_176_nl});
  assign partition_pivot_or_28_nl = (~(swap_equal_tmp_211 | swap_equal_tmp_149 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_14 | swap_1_equal_tmp_78)) & (fsm_output[8]));
  assign partition_pivot_or_29_nl = (swap_equal_tmp_211 & (~ swap_equal_tmp_149)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_14 & (~ swap_1_equal_tmp_78) & (fsm_output[8]));
  assign partition_pivot_or_177_nl = (swap_equal_tmp_149 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_78 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_14_nl = MUX1HOT_v_32_3_2((arr_rsci_din[479:448]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_28_nl , partition_pivot_or_29_nl
      , partition_pivot_or_177_nl});
  assign partition_pivot_or_26_nl = (~(swap_equal_tmp_209 | swap_equal_tmp_147 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_13 | swap_1_equal_tmp_77)) & (fsm_output[8]));
  assign partition_pivot_or_27_nl = (swap_equal_tmp_209 & (~ swap_equal_tmp_147)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_13 & (~ swap_1_equal_tmp_77) & (fsm_output[8]));
  assign partition_pivot_or_178_nl = (swap_equal_tmp_147 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_77 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_13_nl = MUX1HOT_v_32_3_2((arr_rsci_din[447:416]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_26_nl , partition_pivot_or_27_nl
      , partition_pivot_or_178_nl});
  assign partition_pivot_or_24_nl = (~(swap_equal_tmp_207 | swap_equal_tmp_145 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_296 | swap_1_equal_tmp_76)) & (fsm_output[8]));
  assign partition_pivot_or_25_nl = (swap_equal_tmp_207 & (~ swap_equal_tmp_145)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_296 & (~ swap_1_equal_tmp_76) &
      (fsm_output[8]));
  assign partition_pivot_or_179_nl = (swap_equal_tmp_145 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_76 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_12_nl = MUX1HOT_v_32_3_2((arr_rsci_din[415:384]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_24_nl , partition_pivot_or_25_nl
      , partition_pivot_or_179_nl});
  assign partition_pivot_or_22_nl = (~(swap_equal_tmp_205 | swap_equal_tmp_143 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_11 | swap_1_equal_tmp_75)) & (fsm_output[8]));
  assign partition_pivot_or_23_nl = (swap_equal_tmp_205 & (~ swap_equal_tmp_143)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_11 & (~ swap_1_equal_tmp_75) & (fsm_output[8]));
  assign partition_pivot_or_180_nl = (swap_equal_tmp_143 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_75 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_11_nl = MUX1HOT_v_32_3_2((arr_rsci_din[383:352]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_22_nl , partition_pivot_or_23_nl
      , partition_pivot_or_180_nl});
  assign partition_pivot_or_20_nl = (~(swap_equal_tmp_203 | swap_equal_tmp_141 |
      (fsm_output[8]))) | ((~(exit_partition_while_sva | swap_1_equal_tmp_74)) &
      (fsm_output[8]));
  assign partition_pivot_or_21_nl = (swap_equal_tmp_203 & (~ swap_equal_tmp_141)
      & (~ (fsm_output[8]))) | (exit_partition_while_sva & (~ swap_1_equal_tmp_74)
      & (fsm_output[8]));
  assign partition_pivot_or_181_nl = (swap_equal_tmp_141 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_74 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_10_nl = MUX1HOT_v_32_3_2((arr_rsci_din[351:320]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_20_nl , partition_pivot_or_21_nl
      , partition_pivot_or_181_nl});
  assign partition_pivot_or_18_nl = (~(swap_equal_tmp_201 | swap_equal_tmp_139 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_295 | swap_1_equal_tmp_73)) & (fsm_output[8]));
  assign partition_pivot_or_19_nl = (swap_equal_tmp_201 & (~ swap_equal_tmp_139)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_295 & (~ swap_1_equal_tmp_73) &
      (fsm_output[8]));
  assign partition_pivot_or_182_nl = (swap_equal_tmp_139 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_73 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_9_nl = MUX1HOT_v_32_3_2((arr_rsci_din[319:288]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_18_nl , partition_pivot_or_19_nl
      , partition_pivot_or_182_nl});
  assign partition_pivot_or_16_nl = (~(swap_equal_tmp_198 | swap_equal_tmp_199 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_293 | swap_1_equal_tmp_294)) & (fsm_output[8]));
  assign partition_pivot_or_17_nl = (swap_equal_tmp_198 & (~ swap_equal_tmp_199)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_293 & (~ swap_1_equal_tmp_294) &
      (fsm_output[8]));
  assign partition_pivot_or_183_nl = (swap_equal_tmp_199 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_294 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_8_nl = MUX1HOT_v_32_3_2((arr_rsci_din[287:256]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_16_nl , partition_pivot_or_17_nl
      , partition_pivot_or_183_nl});
  assign partition_pivot_or_14_nl = (~(swap_equal_tmp_196 | swap_equal_tmp_136 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_7 | swap_1_equal_tmp_71)) & (fsm_output[8]));
  assign partition_pivot_or_15_nl = (swap_equal_tmp_196 & (~ swap_equal_tmp_136)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_7 & (~ swap_1_equal_tmp_71) & (fsm_output[8]));
  assign partition_pivot_or_184_nl = (swap_equal_tmp_136 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_71 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_7_nl = MUX1HOT_v_32_3_2((arr_rsci_din[255:224]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_14_nl , partition_pivot_or_15_nl
      , partition_pivot_or_184_nl});
  assign partition_pivot_or_12_nl = (~(swap_equal_tmp_193 | swap_equal_tmp_194 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_291 | swap_1_equal_tmp_292)) & (fsm_output[8]));
  assign partition_pivot_or_13_nl = (swap_equal_tmp_193 & (~ swap_equal_tmp_194)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_291 & (~ swap_1_equal_tmp_292) &
      (fsm_output[8]));
  assign partition_pivot_or_185_nl = (swap_equal_tmp_194 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_292 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_6_nl = MUX1HOT_v_32_3_2((arr_rsci_din[223:192]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_12_nl , partition_pivot_or_13_nl
      , partition_pivot_or_185_nl});
  assign partition_pivot_or_10_nl = (~(swap_equal_tmp_190 | swap_equal_tmp_191 |
      (fsm_output[8]))) | ((~(swap_1_equal_tmp_5 | swap_1_equal_tmp_290)) & (fsm_output[8]));
  assign partition_pivot_or_11_nl = (swap_equal_tmp_190 & (~ swap_equal_tmp_191)
      & (~ (fsm_output[8]))) | (swap_1_equal_tmp_5 & (~ swap_1_equal_tmp_290) & (fsm_output[8]));
  assign partition_pivot_or_186_nl = (swap_equal_tmp_191 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_290 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_5_nl = MUX1HOT_v_32_3_2((arr_rsci_din[191:160]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_10_nl , partition_pivot_or_11_nl
      , partition_pivot_or_186_nl});
  assign partition_pivot_or_8_nl = (~(swap_equal_tmp_187 | swap_equal_tmp_188 | (fsm_output[8])))
      | ((~(swap_1_equal_tmp_288 | swap_1_equal_tmp_289)) & (fsm_output[8]));
  assign partition_pivot_or_9_nl = (swap_equal_tmp_187 & (~ swap_equal_tmp_188) &
      (~ (fsm_output[8]))) | (swap_1_equal_tmp_288 & (~ swap_1_equal_tmp_289) & (fsm_output[8]));
  assign partition_pivot_or_187_nl = (swap_equal_tmp_188 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_289 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_4_nl = MUX1HOT_v_32_3_2((arr_rsci_din[159:128]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_8_nl , partition_pivot_or_9_nl
      , partition_pivot_or_187_nl});
  assign partition_pivot_or_6_nl = (~(swap_equal_tmp_184 | swap_equal_tmp_185 | (fsm_output[8])))
      | ((~(swap_1_equal_tmp_3 | swap_1_equal_tmp_287)) & (fsm_output[8]));
  assign partition_pivot_or_7_nl = (swap_equal_tmp_184 & (~ swap_equal_tmp_185) &
      (~ (fsm_output[8]))) | (swap_1_equal_tmp_3 & (~ swap_1_equal_tmp_287) & (fsm_output[8]));
  assign partition_pivot_or_188_nl = (swap_equal_tmp_185 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_287 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_3_nl = MUX1HOT_v_32_3_2((arr_rsci_din[127:96]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_6_nl , partition_pivot_or_7_nl
      , partition_pivot_or_188_nl});
  assign partition_pivot_or_4_nl = (~(swap_equal_tmp_181 | swap_equal_tmp_182 | (fsm_output[8])))
      | ((~(swap_1_equal_tmp_285 | swap_1_equal_tmp_286)) & (fsm_output[8]));
  assign partition_pivot_or_5_nl = (swap_equal_tmp_181 & (~ swap_equal_tmp_182) &
      (~ (fsm_output[8]))) | (swap_1_equal_tmp_285 & (~ swap_1_equal_tmp_286) & (fsm_output[8]));
  assign partition_pivot_or_189_nl = (swap_equal_tmp_182 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_286 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_2_nl = MUX1HOT_v_32_3_2((arr_rsci_din[95:64]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_4_nl , partition_pivot_or_5_nl
      , partition_pivot_or_189_nl});
  assign partition_pivot_or_2_nl = (~(swap_equal_tmp_178 | swap_equal_tmp_179 | (fsm_output[8])))
      | ((~(swap_1_equal_tmp_283 | swap_1_equal_tmp_284)) & (fsm_output[8]));
  assign partition_pivot_or_3_nl = (swap_equal_tmp_178 & (~ swap_equal_tmp_179) &
      (~ (fsm_output[8]))) | (swap_1_equal_tmp_283 & (~ swap_1_equal_tmp_284) & (fsm_output[8]));
  assign partition_pivot_or_190_nl = (swap_equal_tmp_179 & (~ (fsm_output[8]))) |
      (swap_1_equal_tmp_284 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_1_nl = MUX1HOT_v_32_3_2((arr_rsci_din[63:32]),
      partition_while_while_1_mux_2, z_out, {partition_pivot_or_2_nl , partition_pivot_or_3_nl
      , partition_pivot_or_190_nl});
  assign partition_pivot_or_191_nl = (~(swap_or_64_tmp_1 | (fsm_output[8]))) | ((~
      swap_1_or_64_tmp_1) & (fsm_output[8]));
  assign partition_pivot_or_nl = ((~ swap_or_tmp_1) & swap_or_64_tmp_1 & (~ (fsm_output[8])))
      | ((~ swap_1_or_tmp_1) & swap_1_or_64_tmp_1 & (fsm_output[8]));
  assign partition_pivot_or_1_nl = (swap_or_tmp_1 & swap_or_64_tmp_1 & (~ (fsm_output[8])))
      | (swap_1_or_tmp_1 & swap_1_or_64_tmp_1 & (fsm_output[8]));
  assign partition_pivot_partition_pivot_mux1h_nl = MUX1HOT_v_32_3_2(z_out, partition_while_while_1_mux_2,
      (arr_rsci_din[31:0]), {partition_pivot_or_191_nl , partition_pivot_or_nl ,
      partition_pivot_or_1_nl});
  assign nl_arr_rsci_dout = {partition_pivot_partition_pivot_mux1h_63_nl , partition_pivot_partition_pivot_mux1h_62_nl
      , partition_pivot_partition_pivot_mux1h_61_nl , partition_pivot_partition_pivot_mux1h_60_nl
      , partition_pivot_partition_pivot_mux1h_59_nl , partition_pivot_partition_pivot_mux1h_58_nl
      , partition_pivot_partition_pivot_mux1h_57_nl , partition_pivot_partition_pivot_mux1h_56_nl
      , partition_pivot_partition_pivot_mux1h_55_nl , partition_pivot_partition_pivot_mux1h_54_nl
      , partition_pivot_partition_pivot_mux1h_53_nl , partition_pivot_partition_pivot_mux1h_52_nl
      , partition_pivot_partition_pivot_mux1h_51_nl , partition_pivot_partition_pivot_mux1h_50_nl
      , partition_pivot_partition_pivot_mux1h_49_nl , partition_pivot_partition_pivot_mux1h_48_nl
      , partition_pivot_partition_pivot_mux1h_47_nl , partition_pivot_partition_pivot_mux1h_46_nl
      , partition_pivot_partition_pivot_mux1h_45_nl , partition_pivot_partition_pivot_mux1h_44_nl
      , partition_pivot_partition_pivot_mux1h_43_nl , partition_pivot_partition_pivot_mux1h_42_nl
      , partition_pivot_partition_pivot_mux1h_41_nl , partition_pivot_partition_pivot_mux1h_40_nl
      , partition_pivot_partition_pivot_mux1h_39_nl , partition_pivot_partition_pivot_mux1h_38_nl
      , partition_pivot_partition_pivot_mux1h_37_nl , partition_pivot_partition_pivot_mux1h_36_nl
      , partition_pivot_partition_pivot_mux1h_35_nl , partition_pivot_partition_pivot_mux1h_34_nl
      , partition_pivot_partition_pivot_mux1h_33_nl , partition_pivot_partition_pivot_mux1h_32_nl
      , partition_pivot_partition_pivot_mux1h_31_nl , partition_pivot_partition_pivot_mux1h_30_nl
      , partition_pivot_partition_pivot_mux1h_29_nl , partition_pivot_partition_pivot_mux1h_28_nl
      , partition_pivot_partition_pivot_mux1h_27_nl , partition_pivot_partition_pivot_mux1h_26_nl
      , partition_pivot_partition_pivot_mux1h_25_nl , partition_pivot_partition_pivot_mux1h_24_nl
      , partition_pivot_partition_pivot_mux1h_23_nl , partition_pivot_partition_pivot_mux1h_22_nl
      , partition_pivot_partition_pivot_mux1h_21_nl , partition_pivot_partition_pivot_mux1h_20_nl
      , partition_pivot_partition_pivot_mux1h_19_nl , partition_pivot_partition_pivot_mux1h_18_nl
      , partition_pivot_partition_pivot_mux1h_17_nl , partition_pivot_partition_pivot_mux1h_16_nl
      , partition_pivot_partition_pivot_mux1h_15_nl , partition_pivot_partition_pivot_mux1h_14_nl
      , partition_pivot_partition_pivot_mux1h_13_nl , partition_pivot_partition_pivot_mux1h_12_nl
      , partition_pivot_partition_pivot_mux1h_11_nl , partition_pivot_partition_pivot_mux1h_10_nl
      , partition_pivot_partition_pivot_mux1h_9_nl , partition_pivot_partition_pivot_mux1h_8_nl
      , partition_pivot_partition_pivot_mux1h_7_nl , partition_pivot_partition_pivot_mux1h_6_nl
      , partition_pivot_partition_pivot_mux1h_5_nl , partition_pivot_partition_pivot_mux1h_4_nl
      , partition_pivot_partition_pivot_mux1h_3_nl , partition_pivot_partition_pivot_mux1h_2_nl
      , partition_pivot_partition_pivot_mux1h_1_nl , partition_pivot_partition_pivot_mux1h_nl};
  wire  nl_quickSort_core_core_fsm_inst_while_C_0_tr0;
  assign nl_quickSort_core_core_fsm_inst_while_C_0_tr0 = ~ while_acc_3_itm_32_1;
  wire[32:0] partition_while_while_aif_acc_nl;
  wire[33:0] nl_partition_while_while_aif_acc_nl;
  wire  nl_quickSort_core_core_fsm_inst_partition_while_while_C_0_tr0;
  assign nl_partition_while_while_aif_acc_nl = conv_s2u_32_33(z_out_1[31:0]) - conv_s2u_32_33(partition_i_lpi_4);
  assign partition_while_while_aif_acc_nl = nl_partition_while_while_aif_acc_nl[32:0];
  assign nl_quickSort_core_core_fsm_inst_partition_while_while_C_0_tr0 = z_out_2_32
      | (readslicef_33_1_32(partition_while_while_aif_acc_nl));
  wire[32:0] partition_while_while_1_aif_acc_nl;
  wire[33:0] nl_partition_while_while_1_aif_acc_nl;
  wire  nl_quickSort_core_core_fsm_inst_partition_while_while_1_C_0_tr0;
  assign nl_partition_while_while_1_aif_acc_nl = conv_s2u_32_33(partition_j_lpi_4)
      - conv_s2u_32_33(z_out_1[31:0]);
  assign partition_while_while_1_aif_acc_nl = nl_partition_while_while_1_aif_acc_nl[32:0];
  assign nl_quickSort_core_core_fsm_inst_partition_while_while_1_C_0_tr0 = (~ z_out_2_32)
      | (readslicef_33_1_32(partition_while_while_1_aif_acc_nl));
  wire  nl_quickSort_core_core_fsm_inst_while_C_3_tr0;
  assign nl_quickSort_core_core_fsm_inst_while_C_3_tr0 = top_1_31_1_sva_1[30];
  mgc_inout_prereg_en_v1 #(.rscid(32'sd1),
  .width(32'sd2048)) arr_rsci (
      .din(arr_rsci_din),
      .ldout(nl_arr_rsci_ldout),
      .dout(nl_arr_rsci_dout[2047:0]),
      .zin(arr_rsc_zin),
      .lzout(arr_rsc_lzout),
      .zout(arr_rsc_zout)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd32)) low_rsci (
      .dat(low_rsc_dat),
      .idat(low_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd32)) high_rsci (
      .dat(high_rsc_dat),
      .idat(high_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) arr_triosy_obj (
      .ld(reg_high_triosy_obj_ld_cse),
      .lz(arr_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) low_triosy_obj (
      .ld(reg_high_triosy_obj_ld_cse),
      .lz(low_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) high_triosy_obj (
      .ld(reg_high_triosy_obj_ld_cse),
      .lz(high_triosy_lz)
    );
  quickSort_core_core_fsm quickSort_core_core_fsm_inst (
      .clk(clk),
      .rst_n(rst_n),
      .fsm_output(fsm_output),
      .while_C_0_tr0(nl_quickSort_core_core_fsm_inst_while_C_0_tr0),
      .partition_while_while_C_0_tr0(nl_quickSort_core_core_fsm_inst_partition_while_while_C_0_tr0),
      .partition_while_while_1_C_0_tr0(nl_quickSort_core_core_fsm_inst_partition_while_while_1_C_0_tr0),
      .partition_while_C_1_tr0(exit_partition_while_sva),
      .while_C_3_tr0(nl_quickSort_core_core_fsm_inst_while_C_3_tr0)
    );
  assign while_and_1_rgt = while_if_and_122_tmp_sva_1 & while_acc_3_cse_32;
  assign stack_and_1_cse = (while_asn_769 | while_asn_773) & (fsm_output[10]);
  assign stack_and_2_cse = (while_asn_765 | while_asn_769) & (fsm_output[10]);
  assign stack_and_3_cse = (while_asn_761 | while_asn_765) & (fsm_output[10]);
  assign stack_and_4_cse = (while_asn_757 | while_asn_761) & (fsm_output[10]);
  assign stack_and_5_cse = (while_asn_753 | while_asn_757) & (fsm_output[10]);
  assign stack_and_6_cse = (while_asn_749 | while_asn_753) & (fsm_output[10]);
  assign stack_and_7_cse = (while_asn_745 | while_asn_749) & (fsm_output[10]);
  assign stack_and_8_cse = (while_asn_741 | while_asn_745) & (fsm_output[10]);
  assign stack_and_9_cse = (while_asn_737 | while_asn_741) & (fsm_output[10]);
  assign stack_and_10_cse = (while_asn_733 | while_asn_737) & (fsm_output[10]);
  assign stack_and_11_cse = (while_asn_729 | while_asn_733) & (fsm_output[10]);
  assign stack_and_12_cse = (while_asn_725 | while_asn_729) & (fsm_output[10]);
  assign stack_and_13_cse = (while_asn_721 | while_asn_725) & (fsm_output[10]);
  assign stack_and_14_cse = (while_asn_717 | while_asn_721) & (fsm_output[10]);
  assign stack_and_15_cse = (while_asn_713 | while_asn_717) & (fsm_output[10]);
  assign stack_and_16_cse = (while_asn_709 | while_asn_713) & (fsm_output[10]);
  assign stack_and_17_cse = (while_asn_705 | while_asn_709) & (fsm_output[10]);
  assign stack_and_18_cse = (while_asn_701 | while_asn_705) & (fsm_output[10]);
  assign stack_and_19_cse = (while_asn_697 | while_asn_701) & (fsm_output[10]);
  assign stack_and_20_cse = (while_asn_693 | while_asn_697) & (fsm_output[10]);
  assign stack_and_21_cse = (while_asn_689 | while_asn_693) & (fsm_output[10]);
  assign stack_and_22_cse = (while_asn_685 | while_asn_689) & (fsm_output[10]);
  assign stack_and_23_cse = (while_asn_681 | while_asn_685) & (fsm_output[10]);
  assign stack_and_24_cse = (while_asn_677 | while_asn_681) & (fsm_output[10]);
  assign stack_and_25_cse = (while_asn_673 | while_asn_677) & (fsm_output[10]);
  assign stack_and_26_cse = (while_asn_669 | while_asn_673) & (fsm_output[10]);
  assign stack_and_27_cse = (while_asn_665 | while_asn_669) & (fsm_output[10]);
  assign stack_and_28_cse = (while_asn_661 | while_asn_665) & (fsm_output[10]);
  assign stack_and_29_cse = (while_asn_657 | while_asn_661) & (fsm_output[10]);
  assign stack_and_30_cse = (while_asn_653 | while_asn_657) & (fsm_output[10]);
  assign stack_and_31_cse = (while_asn_649 | while_asn_653) & (fsm_output[10]);
  assign stack_and_32_cse = (while_asn_645 | while_asn_649) & (fsm_output[10]);
  assign stack_and_33_cse = (while_asn_641 | while_asn_645) & (fsm_output[10]);
  assign stack_and_34_cse = (while_asn_637 | while_asn_641) & (fsm_output[10]);
  assign stack_and_35_cse = (while_asn_633 | while_asn_637) & (fsm_output[10]);
  assign stack_and_36_cse = (while_asn_629 | while_asn_633) & (fsm_output[10]);
  assign stack_and_37_cse = (while_asn_625 | while_asn_629) & (fsm_output[10]);
  assign stack_and_38_cse = (while_asn_621 | while_asn_625) & (fsm_output[10]);
  assign stack_and_39_cse = (while_asn_617 | while_asn_621) & (fsm_output[10]);
  assign stack_and_40_cse = (while_asn_613 | while_asn_617) & (fsm_output[10]);
  assign stack_and_41_cse = (while_asn_609 | while_asn_613) & (fsm_output[10]);
  assign stack_and_42_cse = (while_asn_605 | while_asn_609) & (fsm_output[10]);
  assign stack_and_43_cse = (while_asn_601 | while_asn_605) & (fsm_output[10]);
  assign stack_and_44_cse = (while_asn_597 | while_asn_601) & (fsm_output[10]);
  assign stack_and_45_cse = (while_asn_593 | while_asn_597) & (fsm_output[10]);
  assign stack_and_46_cse = (while_asn_589 | while_asn_593) & (fsm_output[10]);
  assign stack_and_47_cse = (while_asn_585 | while_asn_589) & (fsm_output[10]);
  assign stack_and_48_cse = (while_asn_581 | while_asn_585) & (fsm_output[10]);
  assign stack_and_49_cse = (while_asn_577 | while_asn_581) & (fsm_output[10]);
  assign stack_and_50_cse = (while_asn_573 | while_asn_577) & (fsm_output[10]);
  assign stack_and_51_cse = (while_asn_569 | while_asn_573) & (fsm_output[10]);
  assign stack_and_52_cse = (while_asn_565 | while_asn_569) & (fsm_output[10]);
  assign stack_and_53_cse = (while_asn_561 | while_asn_565) & (fsm_output[10]);
  assign stack_and_54_cse = (while_asn_557 | while_asn_561) & (fsm_output[10]);
  assign stack_and_55_cse = (while_asn_553 | while_asn_557) & (fsm_output[10]);
  assign stack_and_56_cse = (while_asn_549 | while_asn_553) & (fsm_output[10]);
  assign stack_and_57_cse = (while_asn_545 | while_asn_549) & (fsm_output[10]);
  assign stack_and_58_cse = (while_asn_541 | while_asn_545) & (fsm_output[10]);
  assign stack_and_59_cse = (while_asn_537 | while_asn_541) & (fsm_output[10]);
  assign stack_and_60_cse = (while_asn_533 | while_asn_537) & (fsm_output[10]);
  assign stack_and_61_cse = (while_asn_529 | while_asn_533) & (fsm_output[10]);
  assign stack_and_62_cse = (while_asn_525 | while_asn_529) & (fsm_output[10]);
  assign stack_and_63_cse = (while_asn_523 | while_asn_525) & (fsm_output[10]);
  assign nand_87_cse = ~(and_dcpl_73 & (~ (fsm_output[10])));
  assign nl_while_if_slc_while_if_while_if_acc_tmp = (top_1_31_1_sva_1[29:0]) + 30'b000000000000000000000000000001;
  assign while_if_slc_while_if_while_if_acc_tmp = nl_while_if_slc_while_if_while_if_acc_tmp[29:0];
  assign swap_equal_tmp_128 = (partition_j_lpi_4[5:0]==6'b111111);
  assign swap_equal_tmp_129 = (partition_j_lpi_4[5:0]==6'b111110);
  assign swap_equal_tmp_130 = (partition_j_lpi_4[5:0]==6'b111101);
  assign swap_equal_tmp_131 = (partition_j_lpi_4[5:0]==6'b111100);
  assign swap_equal_tmp_132 = (partition_j_lpi_4[5:0]==6'b111011);
  assign swap_equal_tmp_133 = (partition_j_lpi_4[5:0]==6'b111010);
  assign swap_equal_tmp_134 = (partition_j_lpi_4[5:0]==6'b111001);
  assign swap_equal_tmp_135 = (partition_j_lpi_4[5:0]==6'b111000);
  assign swap_equal_tmp_136 = (partition_j_lpi_4[5:0]==6'b000111);
  assign swap_equal_tmp_137 = (partition_j_lpi_4[5:0]==6'b110111);
  assign swap_equal_tmp_138 = (partition_j_lpi_4[5:0]==6'b110110);
  assign swap_equal_tmp_139 = (partition_j_lpi_4[5:0]==6'b001001);
  assign swap_equal_tmp_140 = (partition_j_lpi_4[5:0]==6'b110101);
  assign swap_equal_tmp_141 = (partition_j_lpi_4[5:0]==6'b001010);
  assign swap_equal_tmp_142 = (partition_j_lpi_4[5:0]==6'b110100);
  assign swap_equal_tmp_143 = (partition_j_lpi_4[5:0]==6'b001011);
  assign swap_equal_tmp_144 = (partition_j_lpi_4[5:0]==6'b110011);
  assign swap_equal_tmp_145 = (partition_j_lpi_4[5:0]==6'b001100);
  assign swap_equal_tmp_146 = (partition_j_lpi_4[5:0]==6'b110010);
  assign swap_equal_tmp_147 = (partition_j_lpi_4[5:0]==6'b001101);
  assign swap_equal_tmp_148 = (partition_j_lpi_4[5:0]==6'b110001);
  assign swap_equal_tmp_149 = (partition_j_lpi_4[5:0]==6'b001110);
  assign swap_equal_tmp_150 = (partition_j_lpi_4[5:0]==6'b001111);
  assign swap_equal_tmp_151 = (partition_j_lpi_4[5:0]==6'b101111);
  assign swap_equal_tmp_152 = (partition_j_lpi_4[5:0]==6'b101110);
  assign swap_equal_tmp_153 = (partition_j_lpi_4[5:0]==6'b101101);
  assign swap_equal_tmp_154 = (partition_j_lpi_4[5:0]==6'b101100);
  assign swap_equal_tmp_155 = (partition_j_lpi_4[5:0]==6'b010011);
  assign swap_equal_tmp_156 = (partition_j_lpi_4[5:0]==6'b101011);
  assign swap_equal_tmp_157 = (partition_j_lpi_4[5:0]==6'b101010);
  assign swap_equal_tmp_158 = (partition_j_lpi_4[5:0]==6'b010101);
  assign swap_equal_tmp_159 = (partition_j_lpi_4[5:0]==6'b101001);
  assign swap_equal_tmp_160 = (partition_j_lpi_4[5:0]==6'b010110);
  assign swap_equal_tmp_161 = (partition_j_lpi_4[5:0]==6'b010111);
  assign swap_equal_tmp_162 = (partition_j_lpi_4[5:0]==6'b100111);
  assign swap_equal_tmp_163 = (partition_j_lpi_4[5:0]==6'b011000);
  assign swap_equal_tmp_164 = (partition_j_lpi_4[5:0]==6'b100110);
  assign swap_equal_tmp_165 = (partition_j_lpi_4[5:0]==6'b011001);
  assign swap_equal_tmp_166 = (partition_j_lpi_4[5:0]==6'b100101);
  assign swap_equal_tmp_167 = (partition_j_lpi_4[5:0]==6'b011010);
  assign swap_equal_tmp_168 = (partition_j_lpi_4[5:0]==6'b100100);
  assign swap_equal_tmp_169 = (partition_j_lpi_4[5:0]==6'b011011);
  assign swap_equal_tmp_170 = (partition_j_lpi_4[5:0]==6'b100011);
  assign swap_equal_tmp_171 = (partition_j_lpi_4[5:0]==6'b011100);
  assign swap_equal_tmp_172 = (partition_j_lpi_4[5:0]==6'b011101);
  assign swap_equal_tmp_173 = (partition_j_lpi_4[5:0]==6'b100001);
  assign swap_equal_tmp_174 = (partition_j_lpi_4[5:0]==6'b011110);
  assign swap_equal_tmp_175 = (partition_j_lpi_4[5:0]==6'b011111);
  assign swap_1_nor_101_itm_1 = ~((partition_j_lpi_4[3:0]!=4'b0000));
  assign while_if_and_369_tmp_sva_1 = while_if_and_stg_4_0_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5);
  assign swap_1_nor_94_itm_2 = ~((partition_j_lpi_4[4]) | (partition_j_lpi_4[2])
      | (partition_j_lpi_4[1]) | (partition_j_lpi_4[0]));
  assign swap_1_nor_88_itm_2 = ~((partition_j_lpi_4[4]) | (partition_j_lpi_4[3])
      | (partition_j_lpi_4[2]) | (partition_j_lpi_4[0]));
  assign swap_1_nor_86_itm_2 = ~((partition_j_lpi_4[4:0]!=5'b00000));
  assign swap_1_nor_75_itm_2 = ~((partition_j_lpi_4[5]) | (partition_j_lpi_4[3])
      | (partition_j_lpi_4[1]) | (partition_j_lpi_4[0]));
  assign swap_1_nor_73_itm_2 = ~((partition_j_lpi_4[5]) | (partition_j_lpi_4[3])
      | (partition_j_lpi_4[2]) | (partition_j_lpi_4[0]));
  assign swap_1_nor_72_itm_2 = ~((partition_j_lpi_4[5]) | (partition_j_lpi_4[3])
      | (partition_j_lpi_4[2]) | (partition_j_lpi_4[1]));
  assign swap_1_nor_71_itm_2 = ~((partition_j_lpi_4[5]) | (partition_j_lpi_4[3])
      | (partition_j_lpi_4[2]) | (partition_j_lpi_4[1]) | (partition_j_lpi_4[0]));
  assign swap_1_nor_63_itm_2 = ~((partition_j_lpi_4[5]) | (partition_j_lpi_4[4])
      | (partition_j_lpi_4[2]) | (partition_j_lpi_4[1]) | (partition_j_lpi_4[0]));
  assign swap_1_nor_61_itm_2 = ~((partition_j_lpi_4[5]) | (partition_j_lpi_4[4])
      | (partition_j_lpi_4[3]) | (partition_j_lpi_4[0]));
  assign swap_1_nor_60_itm_2 = ~((partition_j_lpi_4[5]) | (partition_j_lpi_4[4])
      | (partition_j_lpi_4[3]) | (partition_j_lpi_4[1]));
  assign swap_1_nor_59_itm_2 = ~((partition_j_lpi_4[5]) | (partition_j_lpi_4[4])
      | (partition_j_lpi_4[3]) | (partition_j_lpi_4[1]) | (partition_j_lpi_4[0]));
  assign swap_1_nor_58_itm_1 = ~((partition_j_lpi_4[5:2]!=4'b0000));
  assign while_if_and_stg_4_31_sva_1 = while_if_and_stg_3_15_sva_1 & (partition_pivot_sva_29_0[4]);
  assign swap_1_nor_57_itm_1 = ~((partition_j_lpi_4[5]) | (partition_j_lpi_4[4])
      | (partition_j_lpi_4[3]) | (partition_j_lpi_4[2]) | (partition_j_lpi_4[0]));
  assign while_if_and_stg_4_0_sva_1 = while_if_and_stg_3_0_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign swap_1_nor_56_itm_1 = ~((partition_j_lpi_4[5:1]!=5'b00000));
  assign while_if_and_stg_3_15_sva_1 = while_if_and_stg_2_7_sva_1 & (partition_pivot_sva_29_0[3]);
  assign low_sva_1 = MUX_v_32_64_2(stack_0_1_sva, stack_2_1_sva, stack_4_1_sva, stack_6_1_sva,
      stack_8_1_sva, stack_10_1_sva, stack_12_1_sva, stack_14_1_sva, stack_16_1_sva,
      stack_18_1_sva, stack_20_1_sva, stack_22_1_sva, stack_24_1_sva, stack_26_1_sva,
      stack_28_1_sva, stack_30_1_sva, stack_32_1_sva, stack_34_1_sva, stack_36_1_sva,
      stack_38_1_sva, stack_40_1_sva, stack_42_1_sva, stack_44_1_sva, stack_46_1_sva,
      stack_48_1_sva, stack_50_1_sva, stack_52_1_sva, stack_54_1_sva, stack_56_1_sva,
      stack_58_1_sva, stack_60_1_sva, stack_62_1_sva, stack_64_1_sva, stack_66_1_sva,
      stack_68_1_sva, stack_70_1_sva, stack_72_1_sva, stack_74_1_sva, stack_76_1_sva,
      stack_78_1_sva, stack_80_1_sva, stack_82_1_sva, stack_84_1_sva, stack_86_1_sva,
      stack_88_1_sva, stack_90_1_sva, stack_92_1_sva, stack_94_1_sva, stack_96_1_sva,
      stack_98_1_sva, stack_100_1_sva, stack_102_1_sva, stack_104_1_sva, stack_106_1_sva,
      stack_108_1_sva, stack_110_1_sva, stack_112_1_sva, stack_114_1_sva, stack_116_1_sva,
      stack_118_1_sva, stack_120_1_sva, stack_122_1_sva, stack_124_1_sva, stack_126_1_sva,
      partition_pivot_sva_29_0[5:0]);
  assign while_if_and_stg_2_7_sva_1 = while_if_and_stg_1_3_sva_1 & (partition_pivot_sva_29_0[2]);
  assign while_if_and_stg_1_3_sva_1 = (partition_pivot_sva_29_0[1:0]==2'b11);
  assign while_if_and_stg_1_0_sva_1 = ~((partition_pivot_sva_29_0[1:0]!=2'b00));
  assign while_if_and_stg_3_0_sva_1 = while_if_and_stg_2_0_sva_1 & (~ (partition_pivot_sva_29_0[3]));
  assign while_if_and_stg_2_0_sva_1 = while_if_and_stg_1_0_sva_1 & (~ (partition_pivot_sva_29_0[2]));
  assign while_if_and_122_tmp_sva_1 = while_if_and_stg_4_31_sva_1 & (partition_pivot_sva_29_0[5]);
  assign nl_while_acc_3_nl = conv_s2u_32_33(low_sva_1) - conv_s2u_32_33(high_sva_1);
  assign while_acc_3_nl = nl_while_acc_3_nl[32:0];
  assign while_acc_3_itm_32_1 = readslicef_33_1_32(while_acc_3_nl);
  assign high_sva_1 = MUX_v_32_64_2(stack_1_1_sva, stack_3_1_sva, stack_5_1_sva,
      stack_7_1_sva, stack_9_1_sva, stack_11_1_sva, stack_13_1_sva, stack_15_1_sva,
      stack_17_1_sva, stack_19_1_sva, stack_21_1_sva, stack_23_1_sva, stack_25_1_sva,
      stack_27_1_sva, stack_29_1_sva, stack_31_1_sva, stack_33_1_sva, stack_35_1_sva,
      stack_37_1_sva, stack_39_1_sva, stack_41_1_sva, stack_43_1_sva, stack_45_1_sva,
      stack_47_1_sva, stack_49_1_sva, stack_51_1_sva, stack_53_1_sva, stack_55_1_sva,
      stack_57_1_sva, stack_59_1_sva, stack_61_1_sva, stack_63_1_sva, stack_65_1_sva,
      stack_67_1_sva, stack_69_1_sva, stack_71_1_sva, stack_73_1_sva, stack_75_1_sva,
      stack_77_1_sva, stack_79_1_sva, stack_81_1_sva, stack_83_1_sva, stack_85_1_sva,
      stack_87_1_sva, stack_89_1_sva, stack_91_1_sva, stack_93_1_sva, stack_95_1_sva,
      stack_97_1_sva, stack_99_1_sva, stack_101_1_sva, stack_103_1_sva, stack_105_1_sva,
      stack_107_1_sva, stack_109_1_sva, stack_111_1_sva, stack_113_1_sva, stack_115_1_sva,
      stack_117_1_sva, stack_119_1_sva, stack_121_1_sva, stack_123_1_sva, stack_125_1_sva,
      stack_127_1_sva, partition_pivot_sva_29_0[5:0]);
  assign swap_equal_tmp_176 = (partition_i_lpi_4[5:0]==6'b111111);
  assign partition_while_while_1_mux_2 = MUX_v_32_64_2((arr_rsci_din[31:0]), (arr_rsci_din[63:32]),
      (arr_rsci_din[95:64]), (arr_rsci_din[127:96]), (arr_rsci_din[159:128]), (arr_rsci_din[191:160]),
      (arr_rsci_din[223:192]), (arr_rsci_din[255:224]), (arr_rsci_din[287:256]),
      (arr_rsci_din[319:288]), (arr_rsci_din[351:320]), (arr_rsci_din[383:352]),
      (arr_rsci_din[415:384]), (arr_rsci_din[447:416]), (arr_rsci_din[479:448]),
      (arr_rsci_din[511:480]), (arr_rsci_din[543:512]), (arr_rsci_din[575:544]),
      (arr_rsci_din[607:576]), (arr_rsci_din[639:608]), (arr_rsci_din[671:640]),
      (arr_rsci_din[703:672]), (arr_rsci_din[735:704]), (arr_rsci_din[767:736]),
      (arr_rsci_din[799:768]), (arr_rsci_din[831:800]), (arr_rsci_din[863:832]),
      (arr_rsci_din[895:864]), (arr_rsci_din[927:896]), (arr_rsci_din[959:928]),
      (arr_rsci_din[991:960]), (arr_rsci_din[1023:992]), (arr_rsci_din[1055:1024]),
      (arr_rsci_din[1087:1056]), (arr_rsci_din[1119:1088]), (arr_rsci_din[1151:1120]),
      (arr_rsci_din[1183:1152]), (arr_rsci_din[1215:1184]), (arr_rsci_din[1247:1216]),
      (arr_rsci_din[1279:1248]), (arr_rsci_din[1311:1280]), (arr_rsci_din[1343:1312]),
      (arr_rsci_din[1375:1344]), (arr_rsci_din[1407:1376]), (arr_rsci_din[1439:1408]),
      (arr_rsci_din[1471:1440]), (arr_rsci_din[1503:1472]), (arr_rsci_din[1535:1504]),
      (arr_rsci_din[1567:1536]), (arr_rsci_din[1599:1568]), (arr_rsci_din[1631:1600]),
      (arr_rsci_din[1663:1632]), (arr_rsci_din[1695:1664]), (arr_rsci_din[1727:1696]),
      (arr_rsci_din[1759:1728]), (arr_rsci_din[1791:1760]), (arr_rsci_din[1823:1792]),
      (arr_rsci_din[1855:1824]), (arr_rsci_din[1887:1856]), (arr_rsci_din[1919:1888]),
      (arr_rsci_din[1951:1920]), (arr_rsci_din[1983:1952]), (arr_rsci_din[2015:1984]),
      (arr_rsci_din[2047:2016]), partition_j_lpi_4[5:0]);
  assign swap_or_64_tmp_1 = swap_equal_tmp_179 | swap_equal_tmp_182 | swap_equal_tmp_185
      | swap_equal_tmp_188 | swap_equal_tmp_191 | swap_equal_tmp_194 | swap_equal_tmp_136
      | swap_equal_tmp_199 | swap_equal_tmp_139 | swap_equal_tmp_141 | swap_equal_tmp_143
      | swap_equal_tmp_145 | swap_equal_tmp_147 | swap_equal_tmp_149 | swap_equal_tmp_150
      | swap_equal_tmp_217 | swap_equal_tmp_220 | swap_equal_tmp_223 | swap_equal_tmp_155
      | swap_equal_tmp_228 | swap_equal_tmp_158 | swap_equal_tmp_160 | swap_equal_tmp_161
      | swap_equal_tmp_163 | swap_equal_tmp_165 | swap_equal_tmp_167 | swap_equal_tmp_169
      | swap_equal_tmp_171 | swap_equal_tmp_172 | swap_equal_tmp_174 | swap_equal_tmp_175
      | swap_equal_tmp_252 | swap_equal_tmp_173 | swap_equal_tmp_247 | swap_equal_tmp_170
      | swap_equal_tmp_168 | swap_equal_tmp_166 | swap_equal_tmp_164 | swap_equal_tmp_162
      | swap_equal_tmp_234 | swap_equal_tmp_159 | swap_equal_tmp_157 | swap_equal_tmp_156
      | swap_equal_tmp_154 | swap_equal_tmp_153 | swap_equal_tmp_152 | swap_equal_tmp_151
      | swap_equal_tmp_213 | swap_equal_tmp_148 | swap_equal_tmp_146 | swap_equal_tmp_144
      | swap_equal_tmp_142 | swap_equal_tmp_140 | swap_equal_tmp_138 | swap_equal_tmp_137
      | swap_equal_tmp_135 | swap_equal_tmp_134 | swap_equal_tmp_133 | swap_equal_tmp_132
      | swap_equal_tmp_131 | swap_equal_tmp_130 | swap_equal_tmp_129 | swap_equal_tmp_128;
  assign swap_or_tmp_1 = swap_equal_tmp_178 | swap_equal_tmp_181 | swap_equal_tmp_184
      | swap_equal_tmp_187 | swap_equal_tmp_190 | swap_equal_tmp_193 | swap_equal_tmp_196
      | swap_equal_tmp_198 | swap_equal_tmp_201 | swap_equal_tmp_203 | swap_equal_tmp_205
      | swap_equal_tmp_207 | swap_equal_tmp_209 | swap_equal_tmp_211 | swap_equal_tmp_214
      | swap_equal_tmp_216 | swap_equal_tmp_219 | swap_equal_tmp_222 | swap_equal_tmp_225
      | swap_equal_tmp_227 | swap_equal_tmp_230 | swap_equal_tmp_232 | swap_equal_tmp_235
      | swap_equal_tmp_237 | swap_equal_tmp_239 | swap_equal_tmp_241 | swap_equal_tmp_243
      | swap_equal_tmp_245 | swap_equal_tmp_248 | swap_equal_tmp_250 | swap_equal_tmp_253
      | swap_equal_tmp_251 | swap_equal_tmp_249 | swap_equal_tmp_246 | swap_equal_tmp_244
      | swap_equal_tmp_242 | swap_equal_tmp_240 | swap_equal_tmp_238 | swap_equal_tmp_236
      | swap_equal_tmp_233 | swap_equal_tmp_231 | swap_equal_tmp_229 | swap_equal_tmp_226
      | swap_equal_tmp_224 | swap_equal_tmp_221 | swap_equal_tmp_218 | swap_equal_tmp_215
      | swap_equal_tmp_212 | swap_equal_tmp_210 | swap_equal_tmp_208 | swap_equal_tmp_206
      | swap_equal_tmp_204 | swap_equal_tmp_202 | swap_equal_tmp_200 | swap_equal_tmp_197
      | swap_equal_tmp_195 | swap_equal_tmp_192 | swap_equal_tmp_189 | swap_equal_tmp_186
      | swap_equal_tmp_183 | swap_equal_tmp_180 | swap_equal_tmp_177 | swap_equal_tmp_176;
  assign swap_equal_tmp_177 = (partition_i_lpi_4[5:0]==6'b111110);
  assign swap_equal_tmp_178 = (partition_i_lpi_4[5:0]==6'b000001);
  assign swap_equal_tmp_179 = (partition_j_lpi_4[0]) & swap_1_nor_56_itm_1;
  assign swap_equal_tmp_180 = (partition_i_lpi_4[5:0]==6'b111101);
  assign swap_equal_tmp_181 = (partition_i_lpi_4[5:0]==6'b000010);
  assign swap_equal_tmp_182 = (partition_j_lpi_4[1]) & swap_1_nor_57_itm_1;
  assign swap_equal_tmp_183 = (partition_i_lpi_4[5:0]==6'b111100);
  assign swap_equal_tmp_184 = (partition_i_lpi_4[5:0]==6'b000011);
  assign swap_equal_tmp_185 = (partition_j_lpi_4[1:0]==2'b11) & swap_1_nor_58_itm_1;
  assign swap_equal_tmp_186 = (partition_i_lpi_4[5:0]==6'b111011);
  assign swap_equal_tmp_187 = (partition_i_lpi_4[5:0]==6'b000100);
  assign swap_equal_tmp_188 = (partition_j_lpi_4[2]) & swap_1_nor_59_itm_2;
  assign swap_equal_tmp_189 = (partition_i_lpi_4[5:0]==6'b111010);
  assign swap_equal_tmp_190 = (partition_i_lpi_4[5:0]==6'b000101);
  assign swap_equal_tmp_191 = (partition_j_lpi_4[2]) & (partition_j_lpi_4[0]) & swap_1_nor_60_itm_2;
  assign swap_equal_tmp_192 = (partition_i_lpi_4[5:0]==6'b111001);
  assign swap_equal_tmp_193 = (partition_i_lpi_4[5:0]==6'b000110);
  assign swap_equal_tmp_194 = (partition_j_lpi_4[2:1]==2'b11) & swap_1_nor_61_itm_2;
  assign swap_equal_tmp_195 = (partition_i_lpi_4[5:0]==6'b111000);
  assign swap_equal_tmp_196 = (partition_i_lpi_4[5:0]==6'b000111);
  assign swap_equal_tmp_197 = (partition_i_lpi_4[5:0]==6'b110111);
  assign swap_equal_tmp_198 = (partition_i_lpi_4[5:0]==6'b001000);
  assign swap_equal_tmp_199 = (partition_j_lpi_4[3]) & swap_1_nor_63_itm_2;
  assign swap_equal_tmp_200 = (partition_i_lpi_4[5:0]==6'b110110);
  assign swap_equal_tmp_201 = (partition_i_lpi_4[5:0]==6'b001001);
  assign swap_equal_tmp_202 = (partition_i_lpi_4[5:0]==6'b110101);
  assign swap_equal_tmp_203 = (partition_i_lpi_4[5:0]==6'b001010);
  assign swap_equal_tmp_204 = (partition_i_lpi_4[5:0]==6'b110100);
  assign swap_equal_tmp_205 = (partition_i_lpi_4[5:0]==6'b001011);
  assign swap_equal_tmp_206 = (partition_i_lpi_4[5:0]==6'b110011);
  assign swap_equal_tmp_207 = (partition_i_lpi_4[5:0]==6'b001100);
  assign swap_equal_tmp_208 = (partition_i_lpi_4[5:0]==6'b110010);
  assign swap_equal_tmp_209 = (partition_i_lpi_4[5:0]==6'b001101);
  assign swap_equal_tmp_210 = (partition_i_lpi_4[5:0]==6'b110001);
  assign swap_equal_tmp_211 = (partition_i_lpi_4[5:0]==6'b001110);
  assign swap_equal_tmp_212 = (partition_i_lpi_4[5:0]==6'b110000);
  assign swap_equal_tmp_213 = (partition_j_lpi_4[5:4]==2'b11) & swap_1_nor_101_itm_1;
  assign swap_equal_tmp_214 = (partition_i_lpi_4[5:0]==6'b001111);
  assign swap_equal_tmp_215 = (partition_i_lpi_4[5:0]==6'b101111);
  assign swap_equal_tmp_216 = (partition_i_lpi_4[5:0]==6'b010000);
  assign swap_equal_tmp_217 = (partition_j_lpi_4[4]) & swap_1_nor_71_itm_2;
  assign swap_equal_tmp_218 = (partition_i_lpi_4[5:0]==6'b101110);
  assign swap_equal_tmp_219 = (partition_i_lpi_4[5:0]==6'b010001);
  assign swap_equal_tmp_220 = (partition_j_lpi_4[4]) & (partition_j_lpi_4[0]) & swap_1_nor_72_itm_2;
  assign swap_equal_tmp_221 = (partition_i_lpi_4[5:0]==6'b101101);
  assign swap_equal_tmp_222 = (partition_i_lpi_4[5:0]==6'b010010);
  assign swap_equal_tmp_223 = (partition_j_lpi_4[4]) & (partition_j_lpi_4[1]) & swap_1_nor_73_itm_2;
  assign swap_equal_tmp_224 = (partition_i_lpi_4[5:0]==6'b101100);
  assign swap_equal_tmp_225 = (partition_i_lpi_4[5:0]==6'b010011);
  assign swap_equal_tmp_226 = (partition_i_lpi_4[5:0]==6'b101011);
  assign swap_equal_tmp_227 = (partition_i_lpi_4[5:0]==6'b010100);
  assign swap_equal_tmp_228 = (partition_j_lpi_4[4]) & (partition_j_lpi_4[2]) & swap_1_nor_75_itm_2;
  assign swap_equal_tmp_229 = (partition_i_lpi_4[5:0]==6'b101010);
  assign swap_equal_tmp_230 = (partition_i_lpi_4[5:0]==6'b010101);
  assign swap_equal_tmp_231 = (partition_i_lpi_4[5:0]==6'b101001);
  assign swap_equal_tmp_232 = (partition_i_lpi_4[5:0]==6'b010110);
  assign swap_equal_tmp_233 = (partition_i_lpi_4[5:0]==6'b101000);
  assign swap_equal_tmp_234 = (partition_j_lpi_4[5]) & (partition_j_lpi_4[3]) & swap_1_nor_94_itm_2;
  assign swap_equal_tmp_235 = (partition_i_lpi_4[5:0]==6'b010111);
  assign swap_equal_tmp_236 = (partition_i_lpi_4[5:0]==6'b100111);
  assign swap_equal_tmp_237 = (partition_i_lpi_4[5:0]==6'b011000);
  assign swap_equal_tmp_238 = (partition_i_lpi_4[5:0]==6'b100110);
  assign swap_equal_tmp_239 = (partition_i_lpi_4[5:0]==6'b011001);
  assign swap_equal_tmp_240 = (partition_i_lpi_4[5:0]==6'b100101);
  assign swap_equal_tmp_241 = (partition_i_lpi_4[5:0]==6'b011010);
  assign swap_equal_tmp_242 = (partition_i_lpi_4[5:0]==6'b100100);
  assign swap_equal_tmp_243 = (partition_i_lpi_4[5:0]==6'b011011);
  assign swap_equal_tmp_244 = (partition_i_lpi_4[5:0]==6'b100011);
  assign swap_equal_tmp_245 = (partition_i_lpi_4[5:0]==6'b011100);
  assign swap_equal_tmp_246 = (partition_i_lpi_4[5:0]==6'b100010);
  assign swap_equal_tmp_247 = (partition_j_lpi_4[5]) & (partition_j_lpi_4[1]) & swap_1_nor_88_itm_2;
  assign swap_equal_tmp_248 = (partition_i_lpi_4[5:0]==6'b011101);
  assign swap_equal_tmp_249 = (partition_i_lpi_4[5:0]==6'b100001);
  assign swap_equal_tmp_250 = (partition_i_lpi_4[5:0]==6'b011110);
  assign swap_equal_tmp_251 = (partition_i_lpi_4[5:0]==6'b100000);
  assign swap_equal_tmp_252 = (partition_j_lpi_4[5]) & swap_1_nor_86_itm_2;
  assign swap_equal_tmp_253 = (partition_i_lpi_4[5:0]==6'b011111);
  assign swap_1_or_64_tmp_1 = swap_1_equal_tmp_284 | swap_1_equal_tmp_286 | swap_1_equal_tmp_287
      | swap_1_equal_tmp_289 | swap_1_equal_tmp_290 | swap_1_equal_tmp_292 | swap_1_equal_tmp_71
      | swap_1_equal_tmp_294 | swap_1_equal_tmp_73 | swap_1_equal_tmp_74 | swap_1_equal_tmp_75
      | swap_1_equal_tmp_76 | swap_1_equal_tmp_77 | swap_1_equal_tmp_78 | swap_1_equal_tmp_79
      | swap_1_equal_tmp_299 | swap_1_equal_tmp_300 | swap_1_equal_tmp_301 | swap_1_equal_tmp_83
      | swap_1_equal_tmp_302 | swap_1_equal_tmp_85 | swap_1_equal_tmp_86 | swap_1_equal_tmp_87
      | swap_1_equal_tmp_88 | swap_1_equal_tmp_89 | swap_1_equal_tmp_90 | swap_1_equal_tmp_91
      | swap_1_equal_tmp_92 | swap_1_equal_tmp_93 | swap_1_equal_tmp_94 | swap_1_equal_tmp_95
      | swap_1_equal_tmp_306 | swap_1_equal_tmp_97 | swap_1_equal_tmp_304 | swap_1_equal_tmp_99
      | swap_1_equal_tmp_100 | swap_1_equal_tmp_101 | swap_1_equal_tmp_102 | swap_1_equal_tmp_103
      | swap_1_equal_tmp_303 | swap_1_equal_tmp_105 | swap_1_equal_tmp_106 | swap_1_equal_tmp_107
      | swap_1_equal_tmp_108 | swap_1_equal_tmp_109 | swap_1_equal_tmp_110 | swap_1_equal_tmp_111
      | swap_1_equal_tmp_297 | swap_1_equal_tmp_113 | swap_1_equal_tmp_114 | swap_1_equal_tmp_115
      | swap_1_equal_tmp_116 | swap_1_equal_tmp_117 | swap_1_equal_tmp_118 | swap_1_equal_tmp_119
      | swap_1_equal_tmp_120 | swap_1_equal_tmp_121 | swap_1_equal_tmp_122 | swap_1_equal_tmp_123
      | swap_1_equal_tmp_124 | swap_1_equal_tmp_125 | swap_1_equal_tmp_126 | swap_1_equal_tmp_127;
  assign swap_1_or_tmp_1 = swap_1_equal_tmp_283 | swap_1_equal_tmp_285 | swap_1_equal_tmp_3
      | swap_1_equal_tmp_288 | swap_1_equal_tmp_5 | swap_1_equal_tmp_291 | swap_1_equal_tmp_7
      | swap_1_equal_tmp_293 | swap_1_equal_tmp_295 | exit_partition_while_sva |
      swap_1_equal_tmp_11 | swap_1_equal_tmp_296 | swap_1_equal_tmp_13 | swap_1_equal_tmp_14
      | swap_1_equal_tmp_15 | swap_1_equal_tmp_298 | swap_1_equal_tmp_17 | swap_1_equal_tmp_18
      | swap_1_equal_tmp_19 | swap_1_equal_tmp_20 | swap_1_equal_tmp_21 | swap_1_equal_tmp_22
      | swap_1_equal_tmp_23 | swap_1_equal_tmp_24 | swap_1_equal_tmp_25 | swap_1_equal_tmp_26
      | swap_1_equal_tmp_27 | swap_1_equal_tmp_28 | swap_1_equal_tmp_29 | swap_1_equal_tmp_30
      | swap_1_equal_tmp_31 | swap_1_equal_tmp_305 | swap_1_equal_tmp_33 | swap_1_equal_tmp_34
      | swap_1_equal_tmp_35 | swap_1_equal_tmp_36 | swap_1_equal_tmp_37 | swap_1_equal_tmp_38
      | swap_1_equal_tmp_39 | swap_1_equal_tmp_40 | swap_1_equal_tmp_41 | swap_1_equal_tmp_42
      | swap_1_equal_tmp_43 | swap_1_equal_tmp_44 | swap_1_equal_tmp_45 | swap_1_equal_tmp_46
      | swap_1_equal_tmp_47 | swap_1_equal_tmp_48 | swap_1_equal_tmp_49 | swap_1_equal_tmp_50
      | swap_1_equal_tmp_51 | swap_1_equal_tmp_52 | swap_1_equal_tmp_53 | swap_1_equal_tmp_54
      | swap_1_equal_tmp_55 | swap_1_equal_tmp_56 | swap_1_equal_tmp_57 | swap_1_equal_tmp_58
      | swap_1_equal_tmp_59 | swap_1_equal_tmp_60 | swap_1_equal_tmp_61 | swap_1_equal_tmp_62
      | swap_1_equal_tmp_63;
  assign swap_1_equal_tmp_283 = (low_sva[0]) & swap_1_nor_itm;
  assign swap_1_equal_tmp_284 = (partition_j_lpi_4[0]) & swap_1_nor_56_itm;
  assign swap_1_equal_tmp_285 = (low_sva[1]) & swap_1_nor_1_itm;
  assign swap_1_equal_tmp_286 = (partition_j_lpi_4[1]) & swap_1_nor_57_itm;
  assign swap_1_equal_tmp_287 = (partition_j_lpi_4[1:0]==2'b11) & swap_1_nor_58_itm;
  assign swap_1_equal_tmp_288 = (low_sva[2]) & swap_1_nor_3_itm;
  assign swap_1_equal_tmp_289 = (partition_j_lpi_4[2]) & swap_1_nor_59_itm;
  assign swap_1_equal_tmp_290 = (partition_j_lpi_4[2]) & (partition_j_lpi_4[0]) &
      swap_1_nor_60_itm;
  assign swap_1_equal_tmp_291 = (low_sva[2:1]==2'b11) & swap_1_nor_5_itm;
  assign swap_1_equal_tmp_292 = (partition_j_lpi_4[2:1]==2'b11) & swap_1_nor_61_itm;
  assign swap_1_equal_tmp_293 = (low_sva[3]) & swap_1_nor_7_itm;
  assign swap_1_equal_tmp_294 = (partition_j_lpi_4[3]) & swap_1_nor_63_itm;
  assign swap_1_equal_tmp_295 = (low_sva[3]) & (low_sva[0]) & swap_1_nor_8_itm;
  assign swap_1_equal_tmp_296 = (low_sva[3:2]==2'b11) & swap_1_nor_11_itm;
  assign swap_1_equal_tmp_297 = (partition_j_lpi_4[5:4]==2'b11) & swap_1_nor_101_itm;
  assign swap_1_equal_tmp_298 = (low_sva[4]) & swap_1_nor_15_itm;
  assign swap_1_equal_tmp_299 = (partition_j_lpi_4[4]) & swap_1_nor_71_itm;
  assign swap_1_equal_tmp_300 = (partition_j_lpi_4[4]) & (partition_j_lpi_4[0]) &
      swap_1_nor_72_itm;
  assign swap_1_equal_tmp_301 = (partition_j_lpi_4[4]) & (partition_j_lpi_4[1]) &
      swap_1_nor_73_itm;
  assign swap_1_equal_tmp_302 = (partition_j_lpi_4[4]) & (partition_j_lpi_4[2]) &
      swap_1_nor_75_itm;
  assign swap_1_equal_tmp_303 = (partition_j_lpi_4[5]) & (partition_j_lpi_4[3]) &
      swap_1_nor_94_itm;
  assign swap_1_equal_tmp_304 = (partition_j_lpi_4[5]) & (partition_j_lpi_4[1]) &
      swap_1_nor_88_itm;
  assign swap_1_equal_tmp_305 = (low_sva[5]) & swap_1_nor_30_itm;
  assign swap_1_equal_tmp_306 = (partition_j_lpi_4[5]) & swap_1_nor_86_itm;
  assign while_if_and_stg_4_30_sva_1 = while_if_and_stg_3_14_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_1_sva_1 = while_if_and_stg_3_1_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_29_sva_1 = while_if_and_stg_3_13_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_2_sva_1 = while_if_and_stg_3_2_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_28_sva_1 = while_if_and_stg_3_12_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_3_sva_1 = while_if_and_stg_3_3_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_27_sva_1 = while_if_and_stg_3_11_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_4_sva_1 = while_if_and_stg_3_4_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_26_sva_1 = while_if_and_stg_3_10_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_5_sva_1 = while_if_and_stg_3_5_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_25_sva_1 = while_if_and_stg_3_9_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_6_sva_1 = while_if_and_stg_3_6_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_24_sva_1 = while_if_and_stg_3_8_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_7_sva_1 = while_if_and_stg_3_7_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_23_sva_1 = while_if_and_stg_3_7_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_8_sva_1 = while_if_and_stg_3_8_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_22_sva_1 = while_if_and_stg_3_6_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_9_sva_1 = while_if_and_stg_3_9_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_21_sva_1 = while_if_and_stg_3_5_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_10_sva_1 = while_if_and_stg_3_10_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_20_sva_1 = while_if_and_stg_3_4_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_11_sva_1 = while_if_and_stg_3_11_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_19_sva_1 = while_if_and_stg_3_3_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_12_sva_1 = while_if_and_stg_3_12_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_18_sva_1 = while_if_and_stg_3_2_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_13_sva_1 = while_if_and_stg_3_13_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_17_sva_1 = while_if_and_stg_3_1_sva_1 & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_14_sva_1 = while_if_and_stg_3_14_sva_1 & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_4_16_sva_1 = swap_1_nor_5_itm & (partition_pivot_sva_29_0[4]);
  assign while_if_and_stg_4_15_sva_1 = swap_1_nor_56_itm & (~ (partition_pivot_sva_29_0[4]));
  assign while_if_and_stg_3_1_sva_1 = while_if_and_stg_2_1_sva_1 & (~ (partition_pivot_sva_29_0[3]));
  assign while_if_and_stg_3_2_sva_1 = while_if_and_stg_2_2_sva_1 & (~ (partition_pivot_sva_29_0[3]));
  assign while_if_and_stg_3_3_sva_1 = while_if_and_stg_2_3_sva_1 & (~ (partition_pivot_sva_29_0[3]));
  assign while_if_and_stg_3_4_sva_1 = while_if_and_stg_2_4_sva_1 & (~ (partition_pivot_sva_29_0[3]));
  assign while_if_and_stg_3_5_sva_1 = while_if_and_stg_2_5_sva_1 & (~ (partition_pivot_sva_29_0[3]));
  assign while_if_and_stg_3_6_sva_1 = while_if_and_stg_2_6_sva_1 & (~ (partition_pivot_sva_29_0[3]));
  assign while_if_and_stg_3_7_sva_1 = swap_1_nor_30_itm & (~ (partition_pivot_sva_29_0[3]));
  assign while_if_and_stg_3_8_sva_1 = swap_1_nor_3_itm & (partition_pivot_sva_29_0[3]);
  assign while_if_and_stg_3_9_sva_1 = while_if_and_stg_2_1_sva_1 & (partition_pivot_sva_29_0[3]);
  assign while_if_and_stg_3_10_sva_1 = while_if_and_stg_2_2_sva_1 & (partition_pivot_sva_29_0[3]);
  assign while_if_and_stg_3_11_sva_1 = while_if_and_stg_2_3_sva_1 & (partition_pivot_sva_29_0[3]);
  assign while_if_and_stg_3_12_sva_1 = while_if_and_stg_2_4_sva_1 & (partition_pivot_sva_29_0[3]);
  assign while_if_and_stg_3_13_sva_1 = while_if_and_stg_2_5_sva_1 & (partition_pivot_sva_29_0[3]);
  assign while_if_and_stg_3_14_sva_1 = while_if_and_stg_2_6_sva_1 & (partition_pivot_sva_29_0[3]);
  assign while_if_and_stg_2_1_sva_1 = while_if_and_stg_1_1_sva_1 & (~ (partition_pivot_sva_29_0[2]));
  assign while_if_and_stg_2_2_sva_1 = while_if_and_stg_1_2_sva_1 & (~ (partition_pivot_sva_29_0[2]));
  assign while_if_and_stg_2_3_sva_1 = swap_1_nor_15_itm & (~ (partition_pivot_sva_29_0[2]));
  assign while_if_and_stg_2_4_sva_1 = swap_1_nor_11_itm & (partition_pivot_sva_29_0[2]);
  assign while_if_and_stg_2_5_sva_1 = while_if_and_stg_1_1_sva_1 & (partition_pivot_sva_29_0[2]);
  assign while_if_and_stg_2_6_sva_1 = while_if_and_stg_1_2_sva_1 & (partition_pivot_sva_29_0[2]);
  assign while_if_and_stg_1_1_sva_1 = (partition_pivot_sva_29_0[1:0]==2'b01);
  assign while_if_and_stg_1_2_sva_1 = (partition_pivot_sva_29_0[1:0]==2'b10);
  assign while_asn_523 = swap_1_nor_1_itm & while_acc_3_cse_32;
  assign while_asn_525 = while_if_and_stg_4_30_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_529 = while_if_and_stg_4_29_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_533 = while_if_and_stg_4_28_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_537 = while_if_and_stg_4_27_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_541 = while_if_and_stg_4_26_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_545 = while_if_and_stg_4_25_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_549 = while_if_and_stg_4_24_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_553 = while_if_and_stg_4_23_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_557 = while_if_and_stg_4_22_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_561 = while_if_and_stg_4_21_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_565 = while_if_and_stg_4_20_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_569 = while_if_and_stg_4_19_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_573 = while_if_and_stg_4_18_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_577 = while_if_and_stg_4_17_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_581 = while_if_and_stg_4_16_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_585 = while_if_and_stg_4_15_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_589 = while_if_and_stg_4_14_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_593 = while_if_and_stg_4_13_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_597 = while_if_and_stg_4_12_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_601 = while_if_and_stg_4_11_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_605 = while_if_and_stg_4_10_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_609 = while_if_and_stg_4_9_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_613 = while_if_and_stg_4_8_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_617 = while_if_and_stg_4_7_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_621 = while_if_and_stg_4_6_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_625 = while_if_and_stg_4_5_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_629 = while_if_and_stg_4_4_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_633 = while_if_and_stg_4_3_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_637 = while_if_and_stg_4_2_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_641 = while_if_and_stg_4_1_sva_1 & (partition_pivot_sva_29_0[5])
      & while_acc_3_cse_32;
  assign while_asn_645 = swap_1_nor_57_itm & (partition_pivot_sva_29_0[5]) & while_acc_3_cse_32;
  assign while_asn_649 = swap_1_nor_58_itm & while_if_slc_while_if_while_if_acc_1_psp_sva_5
      & while_acc_3_cse_32;
  assign while_asn_653 = while_if_and_stg_4_30_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_657 = while_if_and_stg_4_29_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_661 = while_if_and_stg_4_28_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_665 = while_if_and_stg_4_27_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_669 = while_if_and_stg_4_26_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_673 = while_if_and_stg_4_25_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_677 = while_if_and_stg_4_24_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_681 = while_if_and_stg_4_23_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_685 = while_if_and_stg_4_22_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_689 = while_if_and_stg_4_21_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_693 = while_if_and_stg_4_20_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_697 = while_if_and_stg_4_19_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_701 = while_if_and_stg_4_18_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_705 = while_if_and_stg_4_17_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_709 = while_if_and_stg_4_16_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_713 = while_if_and_stg_4_15_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_717 = while_if_and_stg_4_14_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_721 = while_if_and_stg_4_13_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_725 = while_if_and_stg_4_12_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_729 = while_if_and_stg_4_11_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_733 = while_if_and_stg_4_10_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_737 = while_if_and_stg_4_9_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_741 = while_if_and_stg_4_8_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_745 = while_if_and_stg_4_7_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_749 = while_if_and_stg_4_6_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_753 = while_if_and_stg_4_5_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_757 = while_if_and_stg_4_4_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_761 = while_if_and_stg_4_3_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_765 = while_if_and_stg_4_2_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_769 = while_if_and_stg_4_1_sva_1 & (~ while_if_slc_while_if_while_if_acc_1_psp_sva_5)
      & while_acc_3_cse_32;
  assign while_asn_773 = swap_1_nor_101_itm & while_acc_3_cse_32;
  assign or_dcpl_1 = (fsm_output[4]) | (fsm_output[2]);
  assign and_dcpl = exit_partition_while_sva & while_acc_3_cse_32;
  assign and_dcpl_73 = ~((fsm_output[0]) | (fsm_output[11]));
  assign or_tmp_613 = and_dcpl_73 & (~((fsm_output[1]) | (fsm_output[10])));
  assign or_tmp_637 = (fsm_output[10]) | (fsm_output[5]);
  assign while_or_193_ssc = (fsm_output[3]) | (fsm_output[6]);
  assign while_or_191_ssc = or_tmp_637 | (fsm_output[9]);
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_0_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( (((while_if_and_369_tmp_sva_1 & while_acc_3_cse_32) | while_and_1_rgt)
        & (~(and_dcpl_73 & (~ (fsm_output[9]))))) | (fsm_output[0]) ) begin
      stack_0_1_sva <= MUX1HOT_v_32_3_2(low_rsci_idat, low_sva, (z_out_1[31:0]),
          {(fsm_output[0]) , and_1186_nl , and_1187_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_2_1_sva <= 32'b00000000000000000000000000000000;
      stack_3_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_1_cse ) begin
      stack_2_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_773);
      stack_3_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_773);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_4_1_sva <= 32'b00000000000000000000000000000000;
      stack_5_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_2_cse ) begin
      stack_4_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_769);
      stack_5_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_769);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_6_1_sva <= 32'b00000000000000000000000000000000;
      stack_7_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_3_cse ) begin
      stack_6_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_765);
      stack_7_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_765);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_8_1_sva <= 32'b00000000000000000000000000000000;
      stack_9_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_4_cse ) begin
      stack_8_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_761);
      stack_9_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_761);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_10_1_sva <= 32'b00000000000000000000000000000000;
      stack_11_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_5_cse ) begin
      stack_10_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_757);
      stack_11_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_757);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_12_1_sva <= 32'b00000000000000000000000000000000;
      stack_13_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_6_cse ) begin
      stack_12_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_753);
      stack_13_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_753);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_14_1_sva <= 32'b00000000000000000000000000000000;
      stack_15_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_7_cse ) begin
      stack_14_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_749);
      stack_15_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_749);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_16_1_sva <= 32'b00000000000000000000000000000000;
      stack_17_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_8_cse ) begin
      stack_16_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_745);
      stack_17_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_745);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_18_1_sva <= 32'b00000000000000000000000000000000;
      stack_19_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_9_cse ) begin
      stack_18_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_741);
      stack_19_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_741);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_20_1_sva <= 32'b00000000000000000000000000000000;
      stack_21_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_10_cse ) begin
      stack_20_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_737);
      stack_21_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_737);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_22_1_sva <= 32'b00000000000000000000000000000000;
      stack_23_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_11_cse ) begin
      stack_22_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_733);
      stack_23_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_733);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_24_1_sva <= 32'b00000000000000000000000000000000;
      stack_25_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_12_cse ) begin
      stack_24_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_729);
      stack_25_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_729);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_26_1_sva <= 32'b00000000000000000000000000000000;
      stack_27_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_13_cse ) begin
      stack_26_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_725);
      stack_27_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_725);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_28_1_sva <= 32'b00000000000000000000000000000000;
      stack_29_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_14_cse ) begin
      stack_28_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_721);
      stack_29_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_721);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_30_1_sva <= 32'b00000000000000000000000000000000;
      stack_31_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_15_cse ) begin
      stack_30_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_717);
      stack_31_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_717);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_32_1_sva <= 32'b00000000000000000000000000000000;
      stack_33_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_16_cse ) begin
      stack_32_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_713);
      stack_33_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_713);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_34_1_sva <= 32'b00000000000000000000000000000000;
      stack_35_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_17_cse ) begin
      stack_34_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_709);
      stack_35_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_709);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_36_1_sva <= 32'b00000000000000000000000000000000;
      stack_37_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_18_cse ) begin
      stack_36_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_705);
      stack_37_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_705);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_38_1_sva <= 32'b00000000000000000000000000000000;
      stack_39_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_19_cse ) begin
      stack_38_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_701);
      stack_39_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_701);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_40_1_sva <= 32'b00000000000000000000000000000000;
      stack_41_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_20_cse ) begin
      stack_40_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_697);
      stack_41_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_697);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_42_1_sva <= 32'b00000000000000000000000000000000;
      stack_43_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_21_cse ) begin
      stack_42_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_693);
      stack_43_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_693);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_44_1_sva <= 32'b00000000000000000000000000000000;
      stack_45_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_22_cse ) begin
      stack_44_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_689);
      stack_45_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_689);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_46_1_sva <= 32'b00000000000000000000000000000000;
      stack_47_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_23_cse ) begin
      stack_46_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_685);
      stack_47_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_685);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_48_1_sva <= 32'b00000000000000000000000000000000;
      stack_49_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_24_cse ) begin
      stack_48_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_681);
      stack_49_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_681);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_50_1_sva <= 32'b00000000000000000000000000000000;
      stack_51_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_25_cse ) begin
      stack_50_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_677);
      stack_51_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_677);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_52_1_sva <= 32'b00000000000000000000000000000000;
      stack_53_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_26_cse ) begin
      stack_52_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_673);
      stack_53_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_673);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_54_1_sva <= 32'b00000000000000000000000000000000;
      stack_55_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_27_cse ) begin
      stack_54_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_669);
      stack_55_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_669);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_56_1_sva <= 32'b00000000000000000000000000000000;
      stack_57_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_28_cse ) begin
      stack_56_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_665);
      stack_57_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_665);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_58_1_sva <= 32'b00000000000000000000000000000000;
      stack_59_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_29_cse ) begin
      stack_58_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_661);
      stack_59_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_661);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_60_1_sva <= 32'b00000000000000000000000000000000;
      stack_61_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_30_cse ) begin
      stack_60_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_657);
      stack_61_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_657);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_62_1_sva <= 32'b00000000000000000000000000000000;
      stack_63_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_31_cse ) begin
      stack_62_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_653);
      stack_63_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_653);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_64_1_sva <= 32'b00000000000000000000000000000000;
      stack_65_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_32_cse ) begin
      stack_64_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_649);
      stack_65_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_649);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_66_1_sva <= 32'b00000000000000000000000000000000;
      stack_67_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_33_cse ) begin
      stack_66_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_645);
      stack_67_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_645);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_68_1_sva <= 32'b00000000000000000000000000000000;
      stack_69_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_34_cse ) begin
      stack_68_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_641);
      stack_69_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_641);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_70_1_sva <= 32'b00000000000000000000000000000000;
      stack_71_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_35_cse ) begin
      stack_70_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_637);
      stack_71_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_637);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_72_1_sva <= 32'b00000000000000000000000000000000;
      stack_73_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_36_cse ) begin
      stack_72_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_633);
      stack_73_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_633);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_74_1_sva <= 32'b00000000000000000000000000000000;
      stack_75_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_37_cse ) begin
      stack_74_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_629);
      stack_75_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_629);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_76_1_sva <= 32'b00000000000000000000000000000000;
      stack_77_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_38_cse ) begin
      stack_76_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_625);
      stack_77_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_625);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_78_1_sva <= 32'b00000000000000000000000000000000;
      stack_79_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_39_cse ) begin
      stack_78_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_621);
      stack_79_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_621);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_80_1_sva <= 32'b00000000000000000000000000000000;
      stack_81_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_40_cse ) begin
      stack_80_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_617);
      stack_81_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_617);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_82_1_sva <= 32'b00000000000000000000000000000000;
      stack_83_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_41_cse ) begin
      stack_82_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_613);
      stack_83_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_613);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_84_1_sva <= 32'b00000000000000000000000000000000;
      stack_85_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_42_cse ) begin
      stack_84_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_609);
      stack_85_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_609);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_86_1_sva <= 32'b00000000000000000000000000000000;
      stack_87_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_43_cse ) begin
      stack_86_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_605);
      stack_87_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_605);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_88_1_sva <= 32'b00000000000000000000000000000000;
      stack_89_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_44_cse ) begin
      stack_88_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_601);
      stack_89_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_601);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_90_1_sva <= 32'b00000000000000000000000000000000;
      stack_91_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_45_cse ) begin
      stack_90_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_597);
      stack_91_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_597);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_92_1_sva <= 32'b00000000000000000000000000000000;
      stack_93_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_46_cse ) begin
      stack_92_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_593);
      stack_93_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_593);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_94_1_sva <= 32'b00000000000000000000000000000000;
      stack_95_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_47_cse ) begin
      stack_94_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_589);
      stack_95_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_589);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_96_1_sva <= 32'b00000000000000000000000000000000;
      stack_97_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_48_cse ) begin
      stack_96_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_585);
      stack_97_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_585);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_98_1_sva <= 32'b00000000000000000000000000000000;
      stack_99_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_49_cse ) begin
      stack_98_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_581);
      stack_99_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_581);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_100_1_sva <= 32'b00000000000000000000000000000000;
      stack_101_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_50_cse ) begin
      stack_100_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_577);
      stack_101_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_577);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_102_1_sva <= 32'b00000000000000000000000000000000;
      stack_103_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_51_cse ) begin
      stack_102_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_573);
      stack_103_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_573);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_104_1_sva <= 32'b00000000000000000000000000000000;
      stack_105_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_52_cse ) begin
      stack_104_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_569);
      stack_105_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_569);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_106_1_sva <= 32'b00000000000000000000000000000000;
      stack_107_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_53_cse ) begin
      stack_106_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_565);
      stack_107_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_565);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_108_1_sva <= 32'b00000000000000000000000000000000;
      stack_109_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_54_cse ) begin
      stack_108_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_561);
      stack_109_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_561);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_110_1_sva <= 32'b00000000000000000000000000000000;
      stack_111_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_55_cse ) begin
      stack_110_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_557);
      stack_111_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_557);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_112_1_sva <= 32'b00000000000000000000000000000000;
      stack_113_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_56_cse ) begin
      stack_112_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_553);
      stack_113_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_553);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_114_1_sva <= 32'b00000000000000000000000000000000;
      stack_115_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_57_cse ) begin
      stack_114_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_549);
      stack_115_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_549);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_116_1_sva <= 32'b00000000000000000000000000000000;
      stack_117_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_58_cse ) begin
      stack_116_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_545);
      stack_117_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_545);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_118_1_sva <= 32'b00000000000000000000000000000000;
      stack_119_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_59_cse ) begin
      stack_118_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_541);
      stack_119_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_541);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_120_1_sva <= 32'b00000000000000000000000000000000;
      stack_121_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_60_cse ) begin
      stack_120_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_537);
      stack_121_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_537);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_122_1_sva <= 32'b00000000000000000000000000000000;
      stack_123_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_61_cse ) begin
      stack_122_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_533);
      stack_123_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_533);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_124_1_sva <= 32'b00000000000000000000000000000000;
      stack_125_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_62_cse ) begin
      stack_124_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_529);
      stack_125_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_529);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_126_1_sva <= 32'b00000000000000000000000000000000;
      stack_127_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( stack_and_63_cse ) begin
      stack_126_1_sva <= MUX_v_32_2_2(low_sva, partition_i_lpi_4, while_asn_525);
      stack_127_1_sva <= MUX_v_32_2_2((z_out_1[31:0]), high_sva, while_asn_525);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      stack_1_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( (((~((~ while_acc_3_cse_32) | exit_partition_while_sva)) | while_asn_773
        | while_asn_523) & nand_87_cse) | (fsm_output[0]) ) begin
      stack_1_1_sva <= MUX1HOT_v_32_3_2(high_rsci_idat, (z_out_1[31:0]), high_sva,
          {(fsm_output[0]) , and_1188_nl , and_1189_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      reg_high_triosy_obj_ld_cse <= 1'b0;
      swap_1_nor_101_itm <= 1'b0;
      swap_1_nor_58_itm <= 1'b0;
      swap_1_nor_57_itm <= 1'b0;
      swap_1_nor_56_itm <= 1'b0;
      swap_1_nor_30_itm <= 1'b0;
      swap_1_nor_15_itm <= 1'b0;
      swap_1_nor_11_itm <= 1'b0;
      swap_1_nor_5_itm <= 1'b0;
      swap_1_nor_3_itm <= 1'b0;
      swap_1_nor_1_itm <= 1'b0;
      exit_partition_while_sva <= 1'b0;
    end
    else begin
      reg_high_triosy_obj_ld_cse <= (top_1_31_1_sva_1[30]) & (fsm_output[10]);
      swap_1_nor_101_itm <= MUX_s_1_2_2(swap_1_nor_101_itm_1, while_if_and_369_tmp_sva_1,
          fsm_output[9]);
      swap_1_nor_58_itm <= MUX_s_1_2_2(swap_1_nor_58_itm_1, while_if_and_stg_4_31_sva_1,
          fsm_output[9]);
      swap_1_nor_57_itm <= MUX_s_1_2_2(swap_1_nor_57_itm_1, while_if_and_stg_4_0_sva_1,
          fsm_output[9]);
      swap_1_nor_56_itm <= MUX_s_1_2_2(swap_1_nor_56_itm_1, while_if_and_stg_3_15_sva_1,
          fsm_output[9]);
      swap_1_nor_30_itm <= MUX_s_1_2_2(swap_1_nor_30_nl, while_if_and_stg_2_7_sva_1,
          fsm_output[9]);
      swap_1_nor_15_itm <= MUX_s_1_2_2(swap_1_nor_15_nl, while_if_and_stg_1_3_sva_1,
          fsm_output[9]);
      swap_1_nor_11_itm <= MUX_s_1_2_2(swap_1_nor_11_nl, while_if_and_stg_1_0_sva_1,
          fsm_output[9]);
      swap_1_nor_5_itm <= MUX_s_1_2_2(swap_1_nor_5_nl, while_if_and_stg_3_0_sva_1,
          fsm_output[9]);
      swap_1_nor_3_itm <= MUX_s_1_2_2(swap_1_nor_3_nl, while_if_and_stg_2_0_sva_1,
          fsm_output[9]);
      swap_1_nor_1_itm <= MUX_s_1_2_2(swap_1_nor_1_nl, while_if_and_122_tmp_sva_1,
          fsm_output[9]);
      exit_partition_while_sva <= MUX1HOT_s_1_3_2((~ (z_out_1[32])), swap_1_swap_1_and_9_nl,
          while_if_while_if_nor_67_nl, {(fsm_output[6]) , (fsm_output[7]) , (fsm_output[9])});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      partition_pivot_sva_31_30 <= 2'b00;
    end
    else if ( ~(or_dcpl_1 | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[7]) |
        (fsm_output[5])) ) begin
      partition_pivot_sva_31_30 <= z_out[31:30];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      partition_pivot_sva_29_0 <= 30'b000000000000000000000000000000;
    end
    else if ( ~((~((fsm_output[7:2]==6'b000000))) | (fsm_output[9])) ) begin
      partition_pivot_sva_29_0 <= MUX_v_30_2_2((z_out[29:0]), and_1160_nl, or_747_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      top_1_31_1_sva_1 <= 31'b0000000000000000000000000000000;
    end
    else if ( ((fsm_output[1]) | (fsm_output[8])) & (while_acc_3_cse_32 | (~ (fsm_output[8])))
        ) begin
      top_1_31_1_sva_1 <= z_out_1[30:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      swap_1_equal_tmp_63 <= 1'b0;
      swap_1_equal_tmp_127 <= 1'b0;
      swap_1_equal_tmp_62 <= 1'b0;
      swap_1_equal_tmp_126 <= 1'b0;
      swap_1_equal_tmp_61 <= 1'b0;
      swap_1_equal_tmp_125 <= 1'b0;
      swap_1_equal_tmp_60 <= 1'b0;
      swap_1_equal_tmp_124 <= 1'b0;
      swap_1_equal_tmp_3 <= 1'b0;
      swap_1_equal_tmp_59 <= 1'b0;
      swap_1_equal_tmp_123 <= 1'b0;
      swap_1_equal_tmp_58 <= 1'b0;
      swap_1_equal_tmp_122 <= 1'b0;
      swap_1_equal_tmp_5 <= 1'b0;
      swap_1_equal_tmp_57 <= 1'b0;
      swap_1_equal_tmp_121 <= 1'b0;
      swap_1_equal_tmp_56 <= 1'b0;
      swap_1_equal_tmp_120 <= 1'b0;
      swap_1_equal_tmp_7 <= 1'b0;
      swap_1_equal_tmp_71 <= 1'b0;
      swap_1_equal_tmp_55 <= 1'b0;
      swap_1_equal_tmp_119 <= 1'b0;
      swap_1_equal_tmp_54 <= 1'b0;
      swap_1_equal_tmp_118 <= 1'b0;
      swap_1_equal_tmp_73 <= 1'b0;
      swap_1_equal_tmp_53 <= 1'b0;
      swap_1_equal_tmp_117 <= 1'b0;
      swap_1_equal_tmp_74 <= 1'b0;
      swap_1_equal_tmp_52 <= 1'b0;
      swap_1_equal_tmp_116 <= 1'b0;
      swap_1_equal_tmp_11 <= 1'b0;
      swap_1_equal_tmp_75 <= 1'b0;
      swap_1_equal_tmp_51 <= 1'b0;
      swap_1_equal_tmp_115 <= 1'b0;
      swap_1_equal_tmp_76 <= 1'b0;
      swap_1_equal_tmp_50 <= 1'b0;
      swap_1_equal_tmp_114 <= 1'b0;
      swap_1_equal_tmp_13 <= 1'b0;
      swap_1_equal_tmp_77 <= 1'b0;
      swap_1_equal_tmp_49 <= 1'b0;
      swap_1_equal_tmp_113 <= 1'b0;
      swap_1_equal_tmp_14 <= 1'b0;
      swap_1_equal_tmp_78 <= 1'b0;
      swap_1_equal_tmp_48 <= 1'b0;
      swap_1_equal_tmp_15 <= 1'b0;
      swap_1_equal_tmp_79 <= 1'b0;
      swap_1_equal_tmp_47 <= 1'b0;
      swap_1_equal_tmp_111 <= 1'b0;
      swap_1_equal_tmp_46 <= 1'b0;
      swap_1_equal_tmp_110 <= 1'b0;
      swap_1_equal_tmp_17 <= 1'b0;
      swap_1_equal_tmp_45 <= 1'b0;
      swap_1_equal_tmp_109 <= 1'b0;
      swap_1_equal_tmp_18 <= 1'b0;
      swap_1_equal_tmp_44 <= 1'b0;
      swap_1_equal_tmp_108 <= 1'b0;
      swap_1_equal_tmp_19 <= 1'b0;
      swap_1_equal_tmp_83 <= 1'b0;
      swap_1_equal_tmp_43 <= 1'b0;
      swap_1_equal_tmp_107 <= 1'b0;
      swap_1_equal_tmp_20 <= 1'b0;
      swap_1_equal_tmp_42 <= 1'b0;
      swap_1_equal_tmp_106 <= 1'b0;
      swap_1_equal_tmp_21 <= 1'b0;
      swap_1_equal_tmp_85 <= 1'b0;
      swap_1_equal_tmp_41 <= 1'b0;
      swap_1_equal_tmp_105 <= 1'b0;
      swap_1_equal_tmp_22 <= 1'b0;
      swap_1_equal_tmp_86 <= 1'b0;
      swap_1_equal_tmp_40 <= 1'b0;
      swap_1_equal_tmp_23 <= 1'b0;
      swap_1_equal_tmp_87 <= 1'b0;
      swap_1_equal_tmp_39 <= 1'b0;
      swap_1_equal_tmp_103 <= 1'b0;
      swap_1_equal_tmp_24 <= 1'b0;
      swap_1_equal_tmp_88 <= 1'b0;
      swap_1_equal_tmp_38 <= 1'b0;
      swap_1_equal_tmp_102 <= 1'b0;
      swap_1_equal_tmp_25 <= 1'b0;
      swap_1_equal_tmp_89 <= 1'b0;
      swap_1_equal_tmp_37 <= 1'b0;
      swap_1_equal_tmp_101 <= 1'b0;
      swap_1_equal_tmp_26 <= 1'b0;
      swap_1_equal_tmp_90 <= 1'b0;
      swap_1_equal_tmp_36 <= 1'b0;
      swap_1_equal_tmp_100 <= 1'b0;
      swap_1_equal_tmp_27 <= 1'b0;
      swap_1_equal_tmp_91 <= 1'b0;
      swap_1_equal_tmp_35 <= 1'b0;
      swap_1_equal_tmp_99 <= 1'b0;
      swap_1_equal_tmp_28 <= 1'b0;
      swap_1_equal_tmp_92 <= 1'b0;
      swap_1_equal_tmp_34 <= 1'b0;
      swap_1_equal_tmp_29 <= 1'b0;
      swap_1_equal_tmp_93 <= 1'b0;
      swap_1_equal_tmp_33 <= 1'b0;
      swap_1_equal_tmp_97 <= 1'b0;
      swap_1_equal_tmp_30 <= 1'b0;
      swap_1_equal_tmp_94 <= 1'b0;
      swap_1_equal_tmp_31 <= 1'b0;
      swap_1_equal_tmp_95 <= 1'b0;
      swap_1_nor_94_itm <= 1'b0;
      swap_1_nor_88_itm <= 1'b0;
      swap_1_nor_86_itm <= 1'b0;
      swap_1_nor_75_itm <= 1'b0;
      swap_1_nor_73_itm <= 1'b0;
      swap_1_nor_72_itm <= 1'b0;
      swap_1_nor_71_itm <= 1'b0;
      swap_1_nor_63_itm <= 1'b0;
      swap_1_nor_61_itm <= 1'b0;
      swap_1_nor_60_itm <= 1'b0;
      swap_1_nor_59_itm <= 1'b0;
      swap_1_nor_8_itm <= 1'b0;
      swap_1_nor_7_itm <= 1'b0;
      swap_1_nor_itm <= 1'b0;
    end
    else if ( and_dcpl ) begin
      swap_1_equal_tmp_63 <= (low_sva[5:0]==6'b111111);
      swap_1_equal_tmp_127 <= swap_equal_tmp_128;
      swap_1_equal_tmp_62 <= (low_sva[5:0]==6'b111110);
      swap_1_equal_tmp_126 <= swap_equal_tmp_129;
      swap_1_equal_tmp_61 <= (low_sva[5:0]==6'b111101);
      swap_1_equal_tmp_125 <= swap_equal_tmp_130;
      swap_1_equal_tmp_60 <= (low_sva[5:0]==6'b111100);
      swap_1_equal_tmp_124 <= swap_equal_tmp_131;
      swap_1_equal_tmp_3 <= (low_sva[5:0]==6'b000011);
      swap_1_equal_tmp_59 <= (low_sva[5:0]==6'b111011);
      swap_1_equal_tmp_123 <= swap_equal_tmp_132;
      swap_1_equal_tmp_58 <= (low_sva[5:0]==6'b111010);
      swap_1_equal_tmp_122 <= swap_equal_tmp_133;
      swap_1_equal_tmp_5 <= (low_sva[5:0]==6'b000101);
      swap_1_equal_tmp_57 <= (low_sva[5:0]==6'b111001);
      swap_1_equal_tmp_121 <= swap_equal_tmp_134;
      swap_1_equal_tmp_56 <= (low_sva[5:0]==6'b111000);
      swap_1_equal_tmp_120 <= swap_equal_tmp_135;
      swap_1_equal_tmp_7 <= (low_sva[5:0]==6'b000111);
      swap_1_equal_tmp_71 <= swap_equal_tmp_136;
      swap_1_equal_tmp_55 <= (low_sva[5:0]==6'b110111);
      swap_1_equal_tmp_119 <= swap_equal_tmp_137;
      swap_1_equal_tmp_54 <= (low_sva[5:0]==6'b110110);
      swap_1_equal_tmp_118 <= swap_equal_tmp_138;
      swap_1_equal_tmp_73 <= swap_equal_tmp_139;
      swap_1_equal_tmp_53 <= (low_sva[5:0]==6'b110101);
      swap_1_equal_tmp_117 <= swap_equal_tmp_140;
      swap_1_equal_tmp_74 <= swap_equal_tmp_141;
      swap_1_equal_tmp_52 <= (low_sva[5:0]==6'b110100);
      swap_1_equal_tmp_116 <= swap_equal_tmp_142;
      swap_1_equal_tmp_11 <= (low_sva[5:0]==6'b001011);
      swap_1_equal_tmp_75 <= swap_equal_tmp_143;
      swap_1_equal_tmp_51 <= (low_sva[5:0]==6'b110011);
      swap_1_equal_tmp_115 <= swap_equal_tmp_144;
      swap_1_equal_tmp_76 <= swap_equal_tmp_145;
      swap_1_equal_tmp_50 <= (low_sva[5:0]==6'b110010);
      swap_1_equal_tmp_114 <= swap_equal_tmp_146;
      swap_1_equal_tmp_13 <= (low_sva[5:0]==6'b001101);
      swap_1_equal_tmp_77 <= swap_equal_tmp_147;
      swap_1_equal_tmp_49 <= (low_sva[5:0]==6'b110001);
      swap_1_equal_tmp_113 <= swap_equal_tmp_148;
      swap_1_equal_tmp_14 <= (low_sva[5:0]==6'b001110);
      swap_1_equal_tmp_78 <= swap_equal_tmp_149;
      swap_1_equal_tmp_48 <= (low_sva[5:0]==6'b110000);
      swap_1_equal_tmp_15 <= (low_sva[5:0]==6'b001111);
      swap_1_equal_tmp_79 <= swap_equal_tmp_150;
      swap_1_equal_tmp_47 <= (low_sva[5:0]==6'b101111);
      swap_1_equal_tmp_111 <= swap_equal_tmp_151;
      swap_1_equal_tmp_46 <= (low_sva[5:0]==6'b101110);
      swap_1_equal_tmp_110 <= swap_equal_tmp_152;
      swap_1_equal_tmp_17 <= (low_sva[5:0]==6'b010001);
      swap_1_equal_tmp_45 <= (low_sva[5:0]==6'b101101);
      swap_1_equal_tmp_109 <= swap_equal_tmp_153;
      swap_1_equal_tmp_18 <= (low_sva[5:0]==6'b010010);
      swap_1_equal_tmp_44 <= (low_sva[5:0]==6'b101100);
      swap_1_equal_tmp_108 <= swap_equal_tmp_154;
      swap_1_equal_tmp_19 <= (low_sva[5:0]==6'b010011);
      swap_1_equal_tmp_83 <= swap_equal_tmp_155;
      swap_1_equal_tmp_43 <= (low_sva[5:0]==6'b101011);
      swap_1_equal_tmp_107 <= swap_equal_tmp_156;
      swap_1_equal_tmp_20 <= (low_sva[5:0]==6'b010100);
      swap_1_equal_tmp_42 <= (low_sva[5:0]==6'b101010);
      swap_1_equal_tmp_106 <= swap_equal_tmp_157;
      swap_1_equal_tmp_21 <= (low_sva[5:0]==6'b010101);
      swap_1_equal_tmp_85 <= swap_equal_tmp_158;
      swap_1_equal_tmp_41 <= (low_sva[5:0]==6'b101001);
      swap_1_equal_tmp_105 <= swap_equal_tmp_159;
      swap_1_equal_tmp_22 <= (low_sva[5:0]==6'b010110);
      swap_1_equal_tmp_86 <= swap_equal_tmp_160;
      swap_1_equal_tmp_40 <= (low_sva[5:0]==6'b101000);
      swap_1_equal_tmp_23 <= (low_sva[5:0]==6'b010111);
      swap_1_equal_tmp_87 <= swap_equal_tmp_161;
      swap_1_equal_tmp_39 <= (low_sva[5:0]==6'b100111);
      swap_1_equal_tmp_103 <= swap_equal_tmp_162;
      swap_1_equal_tmp_24 <= (low_sva[5:0]==6'b011000);
      swap_1_equal_tmp_88 <= swap_equal_tmp_163;
      swap_1_equal_tmp_38 <= (low_sva[5:0]==6'b100110);
      swap_1_equal_tmp_102 <= swap_equal_tmp_164;
      swap_1_equal_tmp_25 <= (low_sva[5:0]==6'b011001);
      swap_1_equal_tmp_89 <= swap_equal_tmp_165;
      swap_1_equal_tmp_37 <= (low_sva[5:0]==6'b100101);
      swap_1_equal_tmp_101 <= swap_equal_tmp_166;
      swap_1_equal_tmp_26 <= (low_sva[5:0]==6'b011010);
      swap_1_equal_tmp_90 <= swap_equal_tmp_167;
      swap_1_equal_tmp_36 <= (low_sva[5:0]==6'b100100);
      swap_1_equal_tmp_100 <= swap_equal_tmp_168;
      swap_1_equal_tmp_27 <= (low_sva[5:0]==6'b011011);
      swap_1_equal_tmp_91 <= swap_equal_tmp_169;
      swap_1_equal_tmp_35 <= (low_sva[5:0]==6'b100011);
      swap_1_equal_tmp_99 <= swap_equal_tmp_170;
      swap_1_equal_tmp_28 <= (low_sva[5:0]==6'b011100);
      swap_1_equal_tmp_92 <= swap_equal_tmp_171;
      swap_1_equal_tmp_34 <= (low_sva[5:0]==6'b100010);
      swap_1_equal_tmp_29 <= (low_sva[5:0]==6'b011101);
      swap_1_equal_tmp_93 <= swap_equal_tmp_172;
      swap_1_equal_tmp_33 <= (low_sva[5:0]==6'b100001);
      swap_1_equal_tmp_97 <= swap_equal_tmp_173;
      swap_1_equal_tmp_30 <= (low_sva[5:0]==6'b011110);
      swap_1_equal_tmp_94 <= swap_equal_tmp_174;
      swap_1_equal_tmp_31 <= (low_sva[5:0]==6'b011111);
      swap_1_equal_tmp_95 <= swap_equal_tmp_175;
      swap_1_nor_94_itm <= swap_1_nor_94_itm_2;
      swap_1_nor_88_itm <= swap_1_nor_88_itm_2;
      swap_1_nor_86_itm <= swap_1_nor_86_itm_2;
      swap_1_nor_75_itm <= swap_1_nor_75_itm_2;
      swap_1_nor_73_itm <= swap_1_nor_73_itm_2;
      swap_1_nor_72_itm <= swap_1_nor_72_itm_2;
      swap_1_nor_71_itm <= swap_1_nor_71_itm_2;
      swap_1_nor_63_itm <= swap_1_nor_63_itm_2;
      swap_1_nor_61_itm <= swap_1_nor_61_itm_2;
      swap_1_nor_60_itm <= swap_1_nor_60_itm_2;
      swap_1_nor_59_itm <= swap_1_nor_59_itm_2;
      swap_1_nor_8_itm <= ~((low_sva[5]) | (low_sva[4]) | (low_sva[2]) | (low_sva[1]));
      swap_1_nor_7_itm <= ~((low_sva[5]) | (low_sva[4]) | (low_sva[2]) | (low_sva[1])
          | (low_sva[0]));
      swap_1_nor_itm <= ~((low_sva[5:1]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      low_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_613 ) begin
      low_sva <= low_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      while_acc_3_cse_32 <= 1'b0;
    end
    else if ( fsm_output[1] ) begin
      while_acc_3_cse_32 <= while_acc_3_itm_32_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      partition_j_lpi_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( nand_87_cse | (fsm_output[1]) | (fsm_output[5]) ) begin
      partition_j_lpi_4 <= MUX_v_32_2_2(high_sva_1, (z_out_1[31:0]), fsm_output[5]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      partition_i_lpi_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( ~(or_dcpl_1 | (fsm_output[7:5]!=3'b000)) ) begin
      partition_i_lpi_4 <= MUX_v_32_2_2(low_sva_1, (z_out_1[31:0]), low_or_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      high_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_613 ) begin
      high_sva <= high_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      while_if_slc_while_if_while_if_acc_1_psp_sva_5 <= 1'b0;
    end
    else if ( ~ (fsm_output[9]) ) begin
      while_if_slc_while_if_while_if_acc_1_psp_sva_5 <= z_out_1[5];
    end
  end
  assign and_1186_nl = (~ while_and_1_rgt) & (fsm_output[9]);
  assign and_1187_nl = while_and_1_rgt & (fsm_output[9]);
  assign and_1188_nl = (~ while_asn_523) & (fsm_output[10]);
  assign and_1189_nl = while_asn_523 & (fsm_output[10]);
  assign swap_1_nor_30_nl = ~((low_sva[4:0]!=5'b00000));
  assign swap_1_nor_15_nl = ~((low_sva[5]) | (low_sva[3]) | (low_sva[2]) | (low_sva[1])
      | (low_sva[0]));
  assign swap_1_nor_11_nl = ~((low_sva[5]) | (low_sva[4]) | (low_sva[1]) | (low_sva[0]));
  assign swap_1_nor_5_nl = ~((low_sva[5]) | (low_sva[4]) | (low_sva[3]) | (low_sva[0]));
  assign swap_1_nor_3_nl = ~((low_sva[5]) | (low_sva[4]) | (low_sva[3]) | (low_sva[1])
      | (low_sva[0]));
  assign swap_1_nor_1_nl = ~((low_sva[5]) | (low_sva[4]) | (low_sva[3]) | (low_sva[2])
      | (low_sva[0]));
  assign swap_1_swap_1_and_9_nl = (low_sva[5:0]==6'b001010);
  assign while_if_while_if_nor_67_nl = ~(while_if_and_369_tmp_sva_1 | while_if_and_122_tmp_sva_1);
  assign mux_nl = MUX_v_30_2_2(while_if_slc_while_if_while_if_acc_tmp, (top_1_31_1_sva_1[29:0]),
      fsm_output[10]);
  assign or_779_nl = (fsm_output[10:8]!=3'b000);
  assign and_1160_nl = MUX_v_30_2_2(30'b000000000000000000000000000000, mux_nl, or_779_nl);
  assign or_747_nl = (fsm_output[0]) | (fsm_output[10]) | (fsm_output[9]) | (fsm_output[8]);
  assign low_or_nl = (fsm_output[3]) | (fsm_output[9]);
  assign while_mux1h_3_nl = MUX1HOT_v_2_4_2((partition_i_lpi_4[31:30]), (partition_j_lpi_4[31:30]),
      (high_sva[31:30]), (low_sva[31:30]), {while_or_193_ssc , while_or_191_ssc ,
      (fsm_output[2]) , (fsm_output[4])});
  assign while_nor_3_nl = ~((fsm_output[1]) | (fsm_output[8]));
  assign while_and_250_nl = MUX_v_2_2_2(2'b00, while_mux1h_3_nl, while_nor_3_nl);
  assign while_mux1h_4_nl = MUX1HOT_v_30_6_2(partition_pivot_sva_29_0, (partition_i_lpi_4[29:0]),
      (partition_j_lpi_4[29:0]), while_if_slc_while_if_while_if_acc_tmp, (high_sva[29:0]),
      (low_sva[29:0]), {(fsm_output[1]) , while_or_193_ssc , while_or_191_ssc , (fsm_output[8])
      , (fsm_output[2]) , (fsm_output[4])});
  assign while_or_196_nl = (~((fsm_output[1]) | (fsm_output[3]) | or_tmp_637 | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[2]) | (fsm_output[4]))) | (fsm_output[6]);
  assign while_mux_1_nl = MUX_v_32_2_2(32'b11111111111111111111111111111110, partition_j_lpi_4,
      fsm_output[6]);
  assign while_nor_5_nl = ~((fsm_output[1]) | or_tmp_637 | (fsm_output[2]));
  assign while_while_while_nand_1_nl = ~(MUX_v_32_2_2(32'b00000000000000000000000000000000,
      while_mux_1_nl, while_nor_5_nl));
  assign nl_acc_nl = conv_s2u_33_34({while_and_250_nl , while_mux1h_4_nl , while_or_196_nl})
      + conv_s2u_33_34({while_while_while_nand_1_nl , 1'b1});
  assign acc_nl = nl_acc_nl[33:0];
  assign z_out_1 = readslicef_34_33_1(acc_nl);
  assign partition_while_while_mux_5_nl = MUX_v_32_2_2((~ z_out), (~ partition_while_while_1_mux_2),
      fsm_output[4]);
  assign nl_acc_1_nl = conv_s2u_33_34({partition_pivot_sva_31_30 , partition_pivot_sva_29_0
      , 1'b1}) + conv_s2u_33_34({partition_while_while_mux_5_nl , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[33:0];
  assign z_out_2_32 = readslicef_34_1_33(acc_1_nl);
  assign or_798_nl = (fsm_output[6]) | (fsm_output[2]);
  assign partition_pivot_mux1h_71_nl = MUX1HOT_v_6_3_2((low_sva_1[5:0]), (partition_i_lpi_4[5:0]),
      (low_sva[5:0]), {(fsm_output[1]) , or_798_nl , (fsm_output[8])});
  assign z_out = MUX_v_32_64_2((arr_rsci_din[31:0]), (arr_rsci_din[63:32]), (arr_rsci_din[95:64]),
      (arr_rsci_din[127:96]), (arr_rsci_din[159:128]), (arr_rsci_din[191:160]), (arr_rsci_din[223:192]),
      (arr_rsci_din[255:224]), (arr_rsci_din[287:256]), (arr_rsci_din[319:288]),
      (arr_rsci_din[351:320]), (arr_rsci_din[383:352]), (arr_rsci_din[415:384]),
      (arr_rsci_din[447:416]), (arr_rsci_din[479:448]), (arr_rsci_din[511:480]),
      (arr_rsci_din[543:512]), (arr_rsci_din[575:544]), (arr_rsci_din[607:576]),
      (arr_rsci_din[639:608]), (arr_rsci_din[671:640]), (arr_rsci_din[703:672]),
      (arr_rsci_din[735:704]), (arr_rsci_din[767:736]), (arr_rsci_din[799:768]),
      (arr_rsci_din[831:800]), (arr_rsci_din[863:832]), (arr_rsci_din[895:864]),
      (arr_rsci_din[927:896]), (arr_rsci_din[959:928]), (arr_rsci_din[991:960]),
      (arr_rsci_din[1023:992]), (arr_rsci_din[1055:1024]), (arr_rsci_din[1087:1056]),
      (arr_rsci_din[1119:1088]), (arr_rsci_din[1151:1120]), (arr_rsci_din[1183:1152]),
      (arr_rsci_din[1215:1184]), (arr_rsci_din[1247:1216]), (arr_rsci_din[1279:1248]),
      (arr_rsci_din[1311:1280]), (arr_rsci_din[1343:1312]), (arr_rsci_din[1375:1344]),
      (arr_rsci_din[1407:1376]), (arr_rsci_din[1439:1408]), (arr_rsci_din[1471:1440]),
      (arr_rsci_din[1503:1472]), (arr_rsci_din[1535:1504]), (arr_rsci_din[1567:1536]),
      (arr_rsci_din[1599:1568]), (arr_rsci_din[1631:1600]), (arr_rsci_din[1663:1632]),
      (arr_rsci_din[1695:1664]), (arr_rsci_din[1727:1696]), (arr_rsci_din[1759:1728]),
      (arr_rsci_din[1791:1760]), (arr_rsci_din[1823:1792]), (arr_rsci_din[1855:1824]),
      (arr_rsci_din[1887:1856]), (arr_rsci_din[1919:1888]), (arr_rsci_din[1951:1920]),
      (arr_rsci_din[1983:1952]), (arr_rsci_din[2015:1984]), (arr_rsci_din[2047:2016]),
      partition_pivot_mux1h_71_nl);

  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_6_2;
    input [29:0] input_5;
    input [29:0] input_4;
    input [29:0] input_3;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [5:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | (input_1 & {30{sel[1]}});
    result = result | (input_2 & {30{sel[2]}});
    result = result | (input_3 & {30{sel[3]}});
    result = result | (input_4 & {30{sel[4]}});
    result = result | (input_5 & {30{sel[5]}});
    MUX1HOT_v_30_6_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | (input_1 & {32{sel[1]}});
    result = result | (input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input  sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_64_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [31:0] input_16;
    input [31:0] input_17;
    input [31:0] input_18;
    input [31:0] input_19;
    input [31:0] input_20;
    input [31:0] input_21;
    input [31:0] input_22;
    input [31:0] input_23;
    input [31:0] input_24;
    input [31:0] input_25;
    input [31:0] input_26;
    input [31:0] input_27;
    input [31:0] input_28;
    input [31:0] input_29;
    input [31:0] input_30;
    input [31:0] input_31;
    input [31:0] input_32;
    input [31:0] input_33;
    input [31:0] input_34;
    input [31:0] input_35;
    input [31:0] input_36;
    input [31:0] input_37;
    input [31:0] input_38;
    input [31:0] input_39;
    input [31:0] input_40;
    input [31:0] input_41;
    input [31:0] input_42;
    input [31:0] input_43;
    input [31:0] input_44;
    input [31:0] input_45;
    input [31:0] input_46;
    input [31:0] input_47;
    input [31:0] input_48;
    input [31:0] input_49;
    input [31:0] input_50;
    input [31:0] input_51;
    input [31:0] input_52;
    input [31:0] input_53;
    input [31:0] input_54;
    input [31:0] input_55;
    input [31:0] input_56;
    input [31:0] input_57;
    input [31:0] input_58;
    input [31:0] input_59;
    input [31:0] input_60;
    input [31:0] input_61;
    input [31:0] input_62;
    input [31:0] input_63;
    input [5:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_32_64_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_34_1_33;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 33;
    readslicef_34_1_33 = tmp[0:0];
  end
  endfunction


  function automatic [32:0] readslicef_34_33_1;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_34_33_1 = tmp[32:0];
  end
  endfunction


  function automatic [32:0] conv_s2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_s2u_32_33 = {vector[31], vector};
  end
  endfunction


  function automatic [33:0] conv_s2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_s2u_33_34 = {vector[32], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    quickSort
// ------------------------------------------------------------------


module quickSort (
  clk, rst_n, arr_rsc_zout, arr_rsc_lzout, arr_rsc_zin, arr_triosy_lz, low_rsc_dat,
      low_triosy_lz, high_rsc_dat, high_triosy_lz
);
  input clk;
  input rst_n;
  output [2047:0] arr_rsc_zout;
  output arr_rsc_lzout;
  input [2047:0] arr_rsc_zin;
  output arr_triosy_lz;
  input [31:0] low_rsc_dat;
  output low_triosy_lz;
  input [31:0] high_rsc_dat;
  output high_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  quickSort_core quickSort_core_inst (
      .clk(clk),
      .rst_n(rst_n),
      .arr_rsc_zout(arr_rsc_zout),
      .arr_rsc_lzout(arr_rsc_lzout),
      .arr_rsc_zin(arr_rsc_zin),
      .arr_triosy_lz(arr_triosy_lz),
      .low_rsc_dat(low_rsc_dat),
      .low_triosy_lz(low_triosy_lz),
      .high_rsc_dat(high_rsc_dat),
      .high_triosy_lz(high_triosy_lz)
    );
endmodule



