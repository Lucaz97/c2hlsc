
//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_inout_prereg_en_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2019 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_inout_prereg_en_v1 (din, ldout, dout, zin, lzout, zout);

    parameter integer rscid = 1;
    parameter integer width = 8;

    output [width-1:0] din;
    input              ldout;
    input  [width-1:0] dout;
    input  [width-1:0] zin;
    output             lzout;
    output [width-1:0] zout;

    wire   [width-1:0] din;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzout = ldout;
    assign din = zin;
    assign zout = dout;

endmodule



//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   lc4976@hansolo.poly.edu
//  Generated date: Tue Apr  9 22:33:57 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    AddRoundKey_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module AddRoundKey_core_core_fsm (
  clk, rst_n, fsm_output, for_C_0_tr0, for_1_for_C_1_tr0, for_1_C_0_tr0
);
  input clk;
  input rst_n;
  output [5:0] fsm_output;
  reg [5:0] fsm_output;
  input for_C_0_tr0;
  input for_1_for_C_1_tr0;
  input for_1_C_0_tr0;


  // FSM State Type Declaration for AddRoundKey_core_core_fsm_1
  parameter
    main_C_0 = 3'd0,
    for_C_0 = 3'd1,
    for_1_for_C_0 = 3'd2,
    for_1_for_C_1 = 3'd3,
    for_1_C_0 = 3'd4,
    main_C_1 = 3'd5;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : AddRoundKey_core_core_fsm_1
    case (state_var)
      for_C_0 : begin
        fsm_output = 6'b000010;
        if ( for_C_0_tr0 ) begin
          state_var_NS = for_1_for_C_0;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      for_1_for_C_0 : begin
        fsm_output = 6'b000100;
        state_var_NS = for_1_for_C_1;
      end
      for_1_for_C_1 : begin
        fsm_output = 6'b001000;
        if ( for_1_for_C_1_tr0 ) begin
          state_var_NS = for_1_C_0;
        end
        else begin
          state_var_NS = for_1_for_C_0;
        end
      end
      for_1_C_0 : begin
        fsm_output = 6'b010000;
        if ( for_1_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_1_for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 6'b100000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 6'b000001;
        state_var_NS = for_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AddRoundKey_core
// ------------------------------------------------------------------


module AddRoundKey_core (
  clk, rst_n, round_rsc_dat, round_triosy_lz, state_rsc_zout, state_rsc_lzout, state_rsc_zin,
      state_triosy_lz, RoundKey_rsc_dat, RoundKey_triosy_lz
);
  input clk;
  input rst_n;
  input [7:0] round_rsc_dat;
  output round_triosy_lz;
  output [127:0] state_rsc_zout;
  output state_rsc_lzout;
  input [127:0] state_rsc_zin;
  output state_triosy_lz;
  input [1415:0] RoundKey_rsc_dat;
  output RoundKey_triosy_lz;


  // Interconnect Declarations
  wire [7:0] round_rsci_idat;
  wire [127:0] state_rsci_din;
  wire [1415:0] RoundKey_rsci_idat;
  wire [5:0] fsm_output;
  wire or_dcpl_1;
  wire or_dcpl_2;
  wire or_dcpl_3;
  wire or_dcpl_4;
  wire or_dcpl_5;
  wire or_dcpl_6;
  wire or_dcpl_7;
  wire or_dcpl_9;
  wire or_dcpl_10;
  wire or_dcpl_12;
  wire or_dcpl_13;
  wire or_dcpl_15;
  wire or_dcpl_16;
  wire or_dcpl_18;
  wire or_dcpl_19;
  wire or_dcpl_21;
  wire or_dcpl_23;
  wire or_dcpl_25;
  wire or_dcpl_27;
  wire or_dcpl_28;
  wire or_dcpl_30;
  wire or_dcpl_32;
  wire or_dcpl_34;
  wire or_dcpl_36;
  wire or_dcpl_37;
  wire or_dcpl_39;
  wire or_dcpl_41;
  wire or_dcpl_43;
  wire or_dcpl_45;
  wire or_dcpl_46;
  wire or_dcpl_63;
  wire or_dcpl_64;
  wire or_dcpl_81;
  wire or_dcpl_82;
  wire or_dcpl_100;
  wire or_dcpl_101;
  wire or_dcpl_118;
  wire or_dcpl_135;
  wire or_dcpl_152;
  wire or_dcpl_169;
  wire or_dcpl_170;
  wire or_dcpl_187;
  wire or_dcpl_204;
  wire or_dcpl_224;
  wire or_dcpl_225;
  wire or_dcpl_226;
  wire or_dcpl_227;
  wire or_dcpl_228;
  wire or_dcpl_229;
  wire or_dcpl_231;
  wire or_dcpl_232;
  wire or_dcpl_234;
  wire or_dcpl_235;
  wire or_dcpl_237;
  wire or_dcpl_238;
  wire or_dcpl_240;
  wire or_dcpl_241;
  wire or_dcpl_243;
  wire or_dcpl_245;
  wire or_dcpl_247;
  wire or_dcpl_249;
  wire or_dcpl_250;
  wire or_dcpl_252;
  wire or_dcpl_254;
  wire or_dcpl_256;
  wire or_dcpl_258;
  wire or_dcpl_259;
  wire or_dcpl_261;
  wire or_dcpl_263;
  wire or_dcpl_265;
  wire or_dcpl_267;
  wire or_dcpl_268;
  wire or_dcpl_285;
  wire or_dcpl_286;
  wire or_dcpl_303;
  wire or_dcpl_304;
  wire or_dcpl_321;
  wire or_dcpl_322;
  wire or_dcpl_339;
  wire or_dcpl_356;
  wire or_dcpl_373;
  wire or_dcpl_390;
  wire or_dcpl_391;
  wire or_dcpl_408;
  wire or_dcpl_425;
  wire or_dcpl_441;
  wire or_dcpl_442;
  wire or_dcpl_444;
  wire or_dcpl_446;
  wire or_dcpl_448;
  wire or_dcpl_449;
  wire or_dcpl_454;
  wire or_dcpl_459;
  reg [7:0] for_slc_i_1_8_7_0_ctmp_sva;
  reg [1:0] i_2_0_sva_1_0;
  reg [1:0] j_2_0_sva_1_0;
  reg reg_RoundKey_triosy_obj_ld_cse;
  wire [7:0] for_1_for_for_1_for_xor_1_cmx_sva_1;
  wire [7:0] z_out;
  wire [8:0] nl_z_out;
  reg [3:0] round_3_0_sva;
  reg [7:0] RoundKey_local_87_sva_1;
  reg [7:0] RoundKey_local_88_sva_1;
  reg [7:0] RoundKey_local_86_sva_1;
  reg [7:0] RoundKey_local_89_sva_1;
  reg [7:0] RoundKey_local_85_sva_1;
  reg [7:0] RoundKey_local_90_sva_1;
  reg [7:0] RoundKey_local_84_sva_1;
  reg [7:0] RoundKey_local_91_sva_1;
  reg [7:0] RoundKey_local_83_sva_1;
  reg [7:0] RoundKey_local_92_sva_1;
  reg [7:0] RoundKey_local_82_sva_1;
  reg [7:0] RoundKey_local_93_sva_1;
  reg [7:0] RoundKey_local_81_sva_1;
  reg [7:0] RoundKey_local_94_sva_1;
  reg [7:0] RoundKey_local_80_sva_1;
  reg [7:0] RoundKey_local_95_sva_1;
  reg [7:0] RoundKey_local_79_sva_1;
  reg [7:0] RoundKey_local_96_sva_1;
  reg [7:0] RoundKey_local_78_sva_1;
  reg [7:0] RoundKey_local_97_sva_1;
  reg [7:0] RoundKey_local_77_sva_1;
  reg [7:0] RoundKey_local_98_sva_1;
  reg [7:0] RoundKey_local_76_sva_1;
  reg [7:0] RoundKey_local_99_sva_1;
  reg [7:0] RoundKey_local_75_sva_1;
  reg [7:0] RoundKey_local_100_sva_1;
  reg [7:0] RoundKey_local_74_sva_1;
  reg [7:0] RoundKey_local_101_sva_1;
  reg [7:0] RoundKey_local_73_sva_1;
  reg [7:0] RoundKey_local_102_sva_1;
  reg [7:0] RoundKey_local_72_sva_1;
  reg [7:0] RoundKey_local_103_sva_1;
  reg [7:0] RoundKey_local_71_sva_1;
  reg [7:0] RoundKey_local_104_sva_1;
  reg [7:0] RoundKey_local_70_sva_1;
  reg [7:0] RoundKey_local_105_sva_1;
  reg [7:0] RoundKey_local_69_sva_1;
  reg [7:0] RoundKey_local_106_sva_1;
  reg [7:0] RoundKey_local_68_sva_1;
  reg [7:0] RoundKey_local_107_sva_1;
  reg [7:0] RoundKey_local_67_sva_1;
  reg [7:0] RoundKey_local_108_sva_1;
  reg [7:0] RoundKey_local_66_sva_1;
  reg [7:0] RoundKey_local_109_sva_1;
  reg [7:0] RoundKey_local_65_sva_1;
  reg [7:0] RoundKey_local_110_sva_1;
  reg [7:0] RoundKey_local_64_sva_1;
  reg [7:0] RoundKey_local_111_sva_1;
  reg [7:0] RoundKey_local_63_sva_1;
  reg [7:0] RoundKey_local_112_sva_1;
  reg [7:0] RoundKey_local_62_sva_1;
  reg [7:0] RoundKey_local_113_sva_1;
  reg [7:0] RoundKey_local_61_sva_1;
  reg [7:0] RoundKey_local_114_sva_1;
  reg [7:0] RoundKey_local_60_sva_1;
  reg [7:0] RoundKey_local_115_sva_1;
  reg [7:0] RoundKey_local_59_sva_1;
  reg [7:0] RoundKey_local_116_sva_1;
  reg [7:0] RoundKey_local_58_sva_1;
  reg [7:0] RoundKey_local_117_sva_1;
  reg [7:0] RoundKey_local_57_sva_1;
  reg [7:0] RoundKey_local_118_sva_1;
  reg [7:0] RoundKey_local_56_sva_1;
  reg [7:0] RoundKey_local_119_sva_1;
  reg [7:0] RoundKey_local_55_sva_1;
  reg [7:0] RoundKey_local_120_sva_1;
  reg [7:0] RoundKey_local_54_sva_1;
  reg [7:0] RoundKey_local_121_sva_1;
  reg [7:0] RoundKey_local_53_sva_1;
  reg [7:0] RoundKey_local_122_sva_1;
  reg [7:0] RoundKey_local_52_sva_1;
  reg [7:0] RoundKey_local_123_sva_1;
  reg [7:0] RoundKey_local_51_sva_1;
  reg [7:0] RoundKey_local_124_sva_1;
  reg [7:0] RoundKey_local_50_sva_1;
  reg [7:0] RoundKey_local_125_sva_1;
  reg [7:0] RoundKey_local_49_sva_1;
  reg [7:0] RoundKey_local_126_sva_1;
  reg [7:0] RoundKey_local_48_sva_1;
  reg [7:0] RoundKey_local_127_sva_1;
  reg [7:0] RoundKey_local_47_sva_1;
  reg [7:0] RoundKey_local_128_sva_1;
  reg [7:0] RoundKey_local_46_sva_1;
  reg [7:0] RoundKey_local_129_sva_1;
  reg [7:0] RoundKey_local_45_sva_1;
  reg [7:0] RoundKey_local_130_sva_1;
  reg [7:0] RoundKey_local_44_sva_1;
  reg [7:0] RoundKey_local_131_sva_1;
  reg [7:0] RoundKey_local_43_sva_1;
  reg [7:0] RoundKey_local_132_sva_1;
  reg [7:0] RoundKey_local_42_sva_1;
  reg [7:0] RoundKey_local_133_sva_1;
  reg [7:0] RoundKey_local_41_sva_1;
  reg [7:0] RoundKey_local_134_sva_1;
  reg [7:0] RoundKey_local_40_sva_1;
  reg [7:0] RoundKey_local_135_sva_1;
  reg [7:0] RoundKey_local_39_sva_1;
  reg [7:0] RoundKey_local_136_sva_1;
  reg [7:0] RoundKey_local_38_sva_1;
  reg [7:0] RoundKey_local_137_sva_1;
  reg [7:0] RoundKey_local_37_sva_1;
  reg [7:0] RoundKey_local_138_sva_1;
  reg [7:0] RoundKey_local_36_sva_1;
  reg [7:0] RoundKey_local_139_sva_1;
  reg [7:0] RoundKey_local_35_sva_1;
  reg [7:0] RoundKey_local_140_sva_1;
  reg [7:0] RoundKey_local_34_sva_1;
  reg [7:0] RoundKey_local_141_sva_1;
  reg [7:0] RoundKey_local_33_sva_1;
  reg [7:0] RoundKey_local_142_sva_1;
  reg [7:0] RoundKey_local_32_sva_1;
  reg [7:0] RoundKey_local_143_sva_1;
  reg [7:0] RoundKey_local_31_sva_1;
  reg [7:0] RoundKey_local_144_sva_1;
  reg [7:0] RoundKey_local_30_sva_1;
  reg [7:0] RoundKey_local_145_sva_1;
  reg [7:0] RoundKey_local_29_sva_1;
  reg [7:0] RoundKey_local_146_sva_1;
  reg [7:0] RoundKey_local_28_sva_1;
  reg [7:0] RoundKey_local_147_sva_1;
  reg [7:0] RoundKey_local_27_sva_1;
  reg [7:0] RoundKey_local_148_sva_1;
  reg [7:0] RoundKey_local_26_sva_1;
  reg [7:0] RoundKey_local_149_sva_1;
  reg [7:0] RoundKey_local_25_sva_1;
  reg [7:0] RoundKey_local_150_sva_1;
  reg [7:0] RoundKey_local_24_sva_1;
  reg [7:0] RoundKey_local_151_sva_1;
  reg [7:0] RoundKey_local_23_sva_1;
  reg [7:0] RoundKey_local_152_sva_1;
  reg [7:0] RoundKey_local_22_sva_1;
  reg [7:0] RoundKey_local_153_sva_1;
  reg [7:0] RoundKey_local_21_sva_1;
  reg [7:0] RoundKey_local_154_sva_1;
  reg [7:0] RoundKey_local_20_sva_1;
  reg [7:0] RoundKey_local_155_sva_1;
  reg [7:0] RoundKey_local_19_sva_1;
  reg [7:0] RoundKey_local_156_sva_1;
  reg [7:0] RoundKey_local_18_sva_1;
  reg [7:0] RoundKey_local_157_sva_1;
  reg [7:0] RoundKey_local_17_sva_1;
  reg [7:0] RoundKey_local_158_sva_1;
  reg [7:0] RoundKey_local_16_sva_1;
  reg [7:0] RoundKey_local_159_sva_1;
  reg [7:0] RoundKey_local_15_sva_1;
  reg [7:0] RoundKey_local_160_sva_1;
  reg [7:0] RoundKey_local_14_sva_1;
  reg [7:0] RoundKey_local_161_sva_1;
  reg [7:0] RoundKey_local_13_sva_1;
  reg [7:0] RoundKey_local_162_sva_1;
  reg [7:0] RoundKey_local_12_sva_1;
  reg [7:0] RoundKey_local_163_sva_1;
  reg [7:0] RoundKey_local_11_sva_1;
  reg [7:0] RoundKey_local_164_sva_1;
  reg [7:0] RoundKey_local_10_sva_1;
  reg [7:0] RoundKey_local_165_sva_1;
  reg [7:0] RoundKey_local_9_sva_1;
  reg [7:0] RoundKey_local_166_sva_1;
  reg [7:0] RoundKey_local_8_sva_1;
  reg [7:0] RoundKey_local_167_sva_1;
  reg [7:0] RoundKey_local_7_sva_1;
  reg [7:0] RoundKey_local_168_sva_1;
  reg [7:0] RoundKey_local_6_sva_1;
  reg [7:0] RoundKey_local_169_sva_1;
  reg [7:0] RoundKey_local_5_sva_1;
  reg [7:0] RoundKey_local_170_sva_1;
  reg [7:0] RoundKey_local_4_sva_1;
  reg [7:0] RoundKey_local_171_sva_1;
  reg [7:0] RoundKey_local_3_sva_1;
  reg [7:0] RoundKey_local_172_sva_1;
  reg [7:0] RoundKey_local_2_sva_1;
  reg [7:0] RoundKey_local_173_sva_1;
  reg [7:0] RoundKey_local_1_sva_1;
  reg [7:0] RoundKey_local_174_sva_1;
  reg [7:0] RoundKey_local_0_sva_1;
  wire [7:0] for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
  wire nor_rgt;
  wire for_acc_itm_4;

  wire[7:0] for_for_mux_nl;
  wire and_372_nl;
  wire[7:0] for_1_for_mux_16_nl;
  wire[7:0] for_1_for_mux_17_nl;
  wire[4:0] for_acc_nl;
  wire[5:0] nl_for_acc_nl;
  wire[5:0] for_for_and_1_nl;
  wire for_nor_2_nl;
  wire[1:0] for_mux1h_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_state_rsci_ldout;
  assign nl_state_rsci_ldout = fsm_output[2];
  wire[7:0] for_1_for_mux_15_nl;
  wire or_466_nl;
  wire[7:0] for_1_for_mux_14_nl;
  wire or_465_nl;
  wire[7:0] for_1_for_mux_13_nl;
  wire or_464_nl;
  wire[7:0] for_1_for_mux_12_nl;
  wire or_463_nl;
  wire[7:0] for_1_for_mux_11_nl;
  wire or_461_nl;
  wire[7:0] for_1_for_mux_10_nl;
  wire or_460_nl;
  wire[7:0] for_1_for_mux_9_nl;
  wire or_459_nl;
  wire[7:0] for_1_for_mux_8_nl;
  wire or_458_nl;
  wire[7:0] for_1_for_mux_7_nl;
  wire or_456_nl;
  wire[7:0] for_1_for_mux_6_nl;
  wire or_455_nl;
  wire[7:0] for_1_for_mux_5_nl;
  wire or_454_nl;
  wire[7:0] for_1_for_mux_4_nl;
  wire or_453_nl;
  wire[7:0] for_1_for_mux_3_nl;
  wire or_450_nl;
  wire[7:0] for_1_for_mux_2_nl;
  wire or_448_nl;
  wire[7:0] for_1_for_mux_1_nl;
  wire or_446_nl;
  wire[7:0] for_1_for_mux_nl;
  wire for_1_for_nor_nl;
  wire [127:0] nl_state_rsci_dout;
  assign or_466_nl = or_dcpl_446 | or_dcpl_459;
  assign for_1_for_mux_15_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[127:120]),
      or_466_nl);
  assign or_465_nl = or_dcpl_444 | or_dcpl_459;
  assign for_1_for_mux_14_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[119:112]),
      or_465_nl);
  assign or_464_nl = or_dcpl_442 | or_dcpl_459;
  assign for_1_for_mux_13_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[111:104]),
      or_464_nl);
  assign or_463_nl = or_dcpl_449 | or_dcpl_459;
  assign for_1_for_mux_12_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[103:96]),
      or_463_nl);
  assign or_461_nl = or_dcpl_446 | or_dcpl_454;
  assign for_1_for_mux_11_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[95:88]),
      or_461_nl);
  assign or_460_nl = or_dcpl_444 | or_dcpl_454;
  assign for_1_for_mux_10_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[87:80]),
      or_460_nl);
  assign or_459_nl = or_dcpl_442 | or_dcpl_454;
  assign for_1_for_mux_9_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[79:72]),
      or_459_nl);
  assign or_458_nl = or_dcpl_449 | or_dcpl_454;
  assign for_1_for_mux_8_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[71:64]),
      or_458_nl);
  assign or_456_nl = or_dcpl_446 | or_dcpl_448;
  assign for_1_for_mux_7_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[63:56]),
      or_456_nl);
  assign or_455_nl = or_dcpl_444 | or_dcpl_448;
  assign for_1_for_mux_6_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[55:48]),
      or_455_nl);
  assign or_454_nl = or_dcpl_442 | or_dcpl_448;
  assign for_1_for_mux_5_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[47:40]),
      or_454_nl);
  assign or_453_nl = or_dcpl_449 | or_dcpl_448;
  assign for_1_for_mux_4_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[39:32]),
      or_453_nl);
  assign or_450_nl = or_dcpl_446 | or_dcpl_441;
  assign for_1_for_mux_3_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[31:24]),
      or_450_nl);
  assign or_448_nl = or_dcpl_444 | or_dcpl_441;
  assign for_1_for_mux_2_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[23:16]),
      or_448_nl);
  assign or_446_nl = or_dcpl_442 | or_dcpl_441;
  assign for_1_for_mux_1_nl = MUX_v_8_2_2(for_1_for_for_1_for_xor_1_cmx_sva_1, (state_rsci_din[15:8]),
      or_446_nl);
  assign for_1_for_nor_nl = ~(((j_2_0_sva_1_0[0]) & (~((i_2_0_sva_1_0!=2'b00) | (j_2_0_sva_1_0[1]))))
      | ((j_2_0_sva_1_0[1]) & (~((i_2_0_sva_1_0!=2'b00) | (j_2_0_sva_1_0[0])))) |
      ((j_2_0_sva_1_0==2'b11) & (i_2_0_sva_1_0==2'b00)) | ((i_2_0_sva_1_0[0]) & (~((i_2_0_sva_1_0[1])
      | (j_2_0_sva_1_0!=2'b00)))) | ((i_2_0_sva_1_0[0]) & (j_2_0_sva_1_0[0]) & (~((i_2_0_sva_1_0[1])
      | (j_2_0_sva_1_0[1])))) | ((i_2_0_sva_1_0[0]) & (j_2_0_sva_1_0[1]) & (~((i_2_0_sva_1_0[1])
      | (j_2_0_sva_1_0[0])))) | ((i_2_0_sva_1_0[0]) & (j_2_0_sva_1_0==2'b11) & (~
      (i_2_0_sva_1_0[1]))) | ((i_2_0_sva_1_0[1]) & (~((i_2_0_sva_1_0[0]) | (j_2_0_sva_1_0!=2'b00))))
      | ((i_2_0_sva_1_0[1]) & (j_2_0_sva_1_0[0]) & (~((i_2_0_sva_1_0[0]) | (j_2_0_sva_1_0[1]))))
      | ((i_2_0_sva_1_0[1]) & (j_2_0_sva_1_0[1]) & (~((i_2_0_sva_1_0[0]) | (j_2_0_sva_1_0[0]))))
      | ((i_2_0_sva_1_0[1]) & (j_2_0_sva_1_0==2'b11) & (~ (i_2_0_sva_1_0[0]))) |
      ((i_2_0_sva_1_0==2'b11) & (j_2_0_sva_1_0==2'b00)) | ((i_2_0_sva_1_0==2'b11)
      & (j_2_0_sva_1_0==2'b01)) | ((i_2_0_sva_1_0==2'b11) & (j_2_0_sva_1_0==2'b10))
      | ((i_2_0_sva_1_0==2'b11) & (j_2_0_sva_1_0==2'b11)));
  assign for_1_for_mux_nl = MUX_v_8_2_2((state_rsci_din[7:0]), for_1_for_for_1_for_xor_1_cmx_sva_1,
      for_1_for_nor_nl);
  assign nl_state_rsci_dout = {for_1_for_mux_15_nl , for_1_for_mux_14_nl , for_1_for_mux_13_nl
      , for_1_for_mux_12_nl , for_1_for_mux_11_nl , for_1_for_mux_10_nl , for_1_for_mux_9_nl
      , for_1_for_mux_8_nl , for_1_for_mux_7_nl , for_1_for_mux_6_nl , for_1_for_mux_5_nl
      , for_1_for_mux_4_nl , for_1_for_mux_3_nl , for_1_for_mux_2_nl , for_1_for_mux_1_nl
      , for_1_for_mux_nl};
  wire  nl_AddRoundKey_core_core_fsm_inst_for_C_0_tr0;
  assign nl_AddRoundKey_core_core_fsm_inst_for_C_0_tr0 = ~ for_acc_itm_4;
  wire  nl_AddRoundKey_core_core_fsm_inst_for_1_for_C_1_tr0;
  assign nl_AddRoundKey_core_core_fsm_inst_for_1_for_C_1_tr0 = z_out[2];
  wire  nl_AddRoundKey_core_core_fsm_inst_for_1_C_0_tr0;
  assign nl_AddRoundKey_core_core_fsm_inst_for_1_C_0_tr0 = z_out[2];
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd8)) round_rsci (
      .dat(round_rsc_dat),
      .idat(round_rsci_idat)
    );
  mgc_inout_prereg_en_v1 #(.rscid(32'sd2),
  .width(32'sd128)) state_rsci (
      .din(state_rsci_din),
      .ldout(nl_state_rsci_ldout),
      .dout(nl_state_rsci_dout[127:0]),
      .zin(state_rsc_zin),
      .lzout(state_rsc_lzout),
      .zout(state_rsc_zout)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd1416)) RoundKey_rsci (
      .dat(RoundKey_rsc_dat),
      .idat(RoundKey_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) round_triosy_obj (
      .ld(reg_RoundKey_triosy_obj_ld_cse),
      .lz(round_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) state_triosy_obj (
      .ld(reg_RoundKey_triosy_obj_ld_cse),
      .lz(state_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) RoundKey_triosy_obj (
      .ld(reg_RoundKey_triosy_obj_ld_cse),
      .lz(RoundKey_triosy_lz)
    );
  AddRoundKey_core_core_fsm AddRoundKey_core_core_fsm_inst (
      .clk(clk),
      .rst_n(rst_n),
      .fsm_output(fsm_output),
      .for_C_0_tr0(nl_AddRoundKey_core_core_fsm_inst_for_C_0_tr0),
      .for_1_for_C_1_tr0(nl_AddRoundKey_core_core_fsm_inst_for_1_for_C_1_tr0),
      .for_1_C_0_tr0(nl_AddRoundKey_core_core_fsm_inst_for_1_C_0_tr0)
    );
  assign nor_rgt = ~((fsm_output[0]) | (fsm_output[5]));
  assign for_slc_i_1_8_7_0_ctmp_sva_mx0w1 = MUX_v_8_176_2((RoundKey_rsci_idat[7:0]),
      (RoundKey_rsci_idat[15:8]), (RoundKey_rsci_idat[23:16]), (RoundKey_rsci_idat[31:24]),
      (RoundKey_rsci_idat[39:32]), (RoundKey_rsci_idat[47:40]), (RoundKey_rsci_idat[55:48]),
      (RoundKey_rsci_idat[63:56]), (RoundKey_rsci_idat[71:64]), (RoundKey_rsci_idat[79:72]),
      (RoundKey_rsci_idat[87:80]), (RoundKey_rsci_idat[95:88]), (RoundKey_rsci_idat[103:96]),
      (RoundKey_rsci_idat[111:104]), (RoundKey_rsci_idat[119:112]), (RoundKey_rsci_idat[127:120]),
      (RoundKey_rsci_idat[135:128]), (RoundKey_rsci_idat[143:136]), (RoundKey_rsci_idat[151:144]),
      (RoundKey_rsci_idat[159:152]), (RoundKey_rsci_idat[167:160]), (RoundKey_rsci_idat[175:168]),
      (RoundKey_rsci_idat[183:176]), (RoundKey_rsci_idat[191:184]), (RoundKey_rsci_idat[199:192]),
      (RoundKey_rsci_idat[207:200]), (RoundKey_rsci_idat[215:208]), (RoundKey_rsci_idat[223:216]),
      (RoundKey_rsci_idat[231:224]), (RoundKey_rsci_idat[239:232]), (RoundKey_rsci_idat[247:240]),
      (RoundKey_rsci_idat[255:248]), (RoundKey_rsci_idat[263:256]), (RoundKey_rsci_idat[271:264]),
      (RoundKey_rsci_idat[279:272]), (RoundKey_rsci_idat[287:280]), (RoundKey_rsci_idat[295:288]),
      (RoundKey_rsci_idat[303:296]), (RoundKey_rsci_idat[311:304]), (RoundKey_rsci_idat[319:312]),
      (RoundKey_rsci_idat[327:320]), (RoundKey_rsci_idat[335:328]), (RoundKey_rsci_idat[343:336]),
      (RoundKey_rsci_idat[351:344]), (RoundKey_rsci_idat[359:352]), (RoundKey_rsci_idat[367:360]),
      (RoundKey_rsci_idat[375:368]), (RoundKey_rsci_idat[383:376]), (RoundKey_rsci_idat[391:384]),
      (RoundKey_rsci_idat[399:392]), (RoundKey_rsci_idat[407:400]), (RoundKey_rsci_idat[415:408]),
      (RoundKey_rsci_idat[423:416]), (RoundKey_rsci_idat[431:424]), (RoundKey_rsci_idat[439:432]),
      (RoundKey_rsci_idat[447:440]), (RoundKey_rsci_idat[455:448]), (RoundKey_rsci_idat[463:456]),
      (RoundKey_rsci_idat[471:464]), (RoundKey_rsci_idat[479:472]), (RoundKey_rsci_idat[487:480]),
      (RoundKey_rsci_idat[495:488]), (RoundKey_rsci_idat[503:496]), (RoundKey_rsci_idat[511:504]),
      (RoundKey_rsci_idat[519:512]), (RoundKey_rsci_idat[527:520]), (RoundKey_rsci_idat[535:528]),
      (RoundKey_rsci_idat[543:536]), (RoundKey_rsci_idat[551:544]), (RoundKey_rsci_idat[559:552]),
      (RoundKey_rsci_idat[567:560]), (RoundKey_rsci_idat[575:568]), (RoundKey_rsci_idat[583:576]),
      (RoundKey_rsci_idat[591:584]), (RoundKey_rsci_idat[599:592]), (RoundKey_rsci_idat[607:600]),
      (RoundKey_rsci_idat[615:608]), (RoundKey_rsci_idat[623:616]), (RoundKey_rsci_idat[631:624]),
      (RoundKey_rsci_idat[639:632]), (RoundKey_rsci_idat[647:640]), (RoundKey_rsci_idat[655:648]),
      (RoundKey_rsci_idat[663:656]), (RoundKey_rsci_idat[671:664]), (RoundKey_rsci_idat[679:672]),
      (RoundKey_rsci_idat[687:680]), (RoundKey_rsci_idat[695:688]), (RoundKey_rsci_idat[703:696]),
      (RoundKey_rsci_idat[711:704]), (RoundKey_rsci_idat[719:712]), (RoundKey_rsci_idat[727:720]),
      (RoundKey_rsci_idat[735:728]), (RoundKey_rsci_idat[743:736]), (RoundKey_rsci_idat[751:744]),
      (RoundKey_rsci_idat[759:752]), (RoundKey_rsci_idat[767:760]), (RoundKey_rsci_idat[775:768]),
      (RoundKey_rsci_idat[783:776]), (RoundKey_rsci_idat[791:784]), (RoundKey_rsci_idat[799:792]),
      (RoundKey_rsci_idat[807:800]), (RoundKey_rsci_idat[815:808]), (RoundKey_rsci_idat[823:816]),
      (RoundKey_rsci_idat[831:824]), (RoundKey_rsci_idat[839:832]), (RoundKey_rsci_idat[847:840]),
      (RoundKey_rsci_idat[855:848]), (RoundKey_rsci_idat[863:856]), (RoundKey_rsci_idat[871:864]),
      (RoundKey_rsci_idat[879:872]), (RoundKey_rsci_idat[887:880]), (RoundKey_rsci_idat[895:888]),
      (RoundKey_rsci_idat[903:896]), (RoundKey_rsci_idat[911:904]), (RoundKey_rsci_idat[919:912]),
      (RoundKey_rsci_idat[927:920]), (RoundKey_rsci_idat[935:928]), (RoundKey_rsci_idat[943:936]),
      (RoundKey_rsci_idat[951:944]), (RoundKey_rsci_idat[959:952]), (RoundKey_rsci_idat[967:960]),
      (RoundKey_rsci_idat[975:968]), (RoundKey_rsci_idat[983:976]), (RoundKey_rsci_idat[991:984]),
      (RoundKey_rsci_idat[999:992]), (RoundKey_rsci_idat[1007:1000]), (RoundKey_rsci_idat[1015:1008]),
      (RoundKey_rsci_idat[1023:1016]), (RoundKey_rsci_idat[1031:1024]), (RoundKey_rsci_idat[1039:1032]),
      (RoundKey_rsci_idat[1047:1040]), (RoundKey_rsci_idat[1055:1048]), (RoundKey_rsci_idat[1063:1056]),
      (RoundKey_rsci_idat[1071:1064]), (RoundKey_rsci_idat[1079:1072]), (RoundKey_rsci_idat[1087:1080]),
      (RoundKey_rsci_idat[1095:1088]), (RoundKey_rsci_idat[1103:1096]), (RoundKey_rsci_idat[1111:1104]),
      (RoundKey_rsci_idat[1119:1112]), (RoundKey_rsci_idat[1127:1120]), (RoundKey_rsci_idat[1135:1128]),
      (RoundKey_rsci_idat[1143:1136]), (RoundKey_rsci_idat[1151:1144]), (RoundKey_rsci_idat[1159:1152]),
      (RoundKey_rsci_idat[1167:1160]), (RoundKey_rsci_idat[1175:1168]), (RoundKey_rsci_idat[1183:1176]),
      (RoundKey_rsci_idat[1191:1184]), (RoundKey_rsci_idat[1199:1192]), (RoundKey_rsci_idat[1207:1200]),
      (RoundKey_rsci_idat[1215:1208]), (RoundKey_rsci_idat[1223:1216]), (RoundKey_rsci_idat[1231:1224]),
      (RoundKey_rsci_idat[1239:1232]), (RoundKey_rsci_idat[1247:1240]), (RoundKey_rsci_idat[1255:1248]),
      (RoundKey_rsci_idat[1263:1256]), (RoundKey_rsci_idat[1271:1264]), (RoundKey_rsci_idat[1279:1272]),
      (RoundKey_rsci_idat[1287:1280]), (RoundKey_rsci_idat[1295:1288]), (RoundKey_rsci_idat[1303:1296]),
      (RoundKey_rsci_idat[1311:1304]), (RoundKey_rsci_idat[1319:1312]), (RoundKey_rsci_idat[1327:1320]),
      (RoundKey_rsci_idat[1335:1328]), (RoundKey_rsci_idat[1343:1336]), (RoundKey_rsci_idat[1351:1344]),
      (RoundKey_rsci_idat[1359:1352]), (RoundKey_rsci_idat[1367:1360]), (RoundKey_rsci_idat[1375:1368]),
      (RoundKey_rsci_idat[1383:1376]), (RoundKey_rsci_idat[1391:1384]), (RoundKey_rsci_idat[1399:1392]),
      (RoundKey_rsci_idat[1407:1400]), for_slc_i_1_8_7_0_ctmp_sva);
  assign for_1_for_mux_16_nl = MUX_v_8_16_2((state_rsci_din[7:0]), (state_rsci_din[15:8]),
      (state_rsci_din[23:16]), (state_rsci_din[31:24]), (state_rsci_din[39:32]),
      (state_rsci_din[47:40]), (state_rsci_din[55:48]), (state_rsci_din[63:56]),
      (state_rsci_din[71:64]), (state_rsci_din[79:72]), (state_rsci_din[87:80]),
      (state_rsci_din[95:88]), (state_rsci_din[103:96]), (state_rsci_din[111:104]),
      (state_rsci_din[119:112]), (state_rsci_din[127:120]), {i_2_0_sva_1_0 , j_2_0_sva_1_0});
  assign for_1_for_mux_17_nl = MUX_v_8_176_2(RoundKey_local_0_sva_1, RoundKey_local_1_sva_1,
      RoundKey_local_2_sva_1, RoundKey_local_3_sva_1, RoundKey_local_4_sva_1, RoundKey_local_5_sva_1,
      RoundKey_local_6_sva_1, RoundKey_local_7_sva_1, RoundKey_local_8_sva_1, RoundKey_local_9_sva_1,
      RoundKey_local_10_sva_1, RoundKey_local_11_sva_1, RoundKey_local_12_sva_1,
      RoundKey_local_13_sva_1, RoundKey_local_14_sva_1, RoundKey_local_15_sva_1,
      RoundKey_local_16_sva_1, RoundKey_local_17_sva_1, RoundKey_local_18_sva_1,
      RoundKey_local_19_sva_1, RoundKey_local_20_sva_1, RoundKey_local_21_sva_1,
      RoundKey_local_22_sva_1, RoundKey_local_23_sva_1, RoundKey_local_24_sva_1,
      RoundKey_local_25_sva_1, RoundKey_local_26_sva_1, RoundKey_local_27_sva_1,
      RoundKey_local_28_sva_1, RoundKey_local_29_sva_1, RoundKey_local_30_sva_1,
      RoundKey_local_31_sva_1, RoundKey_local_32_sva_1, RoundKey_local_33_sva_1,
      RoundKey_local_34_sva_1, RoundKey_local_35_sva_1, RoundKey_local_36_sva_1,
      RoundKey_local_37_sva_1, RoundKey_local_38_sva_1, RoundKey_local_39_sva_1,
      RoundKey_local_40_sva_1, RoundKey_local_41_sva_1, RoundKey_local_42_sva_1,
      RoundKey_local_43_sva_1, RoundKey_local_44_sva_1, RoundKey_local_45_sva_1,
      RoundKey_local_46_sva_1, RoundKey_local_47_sva_1, RoundKey_local_48_sva_1,
      RoundKey_local_49_sva_1, RoundKey_local_50_sva_1, RoundKey_local_51_sva_1,
      RoundKey_local_52_sva_1, RoundKey_local_53_sva_1, RoundKey_local_54_sva_1,
      RoundKey_local_55_sva_1, RoundKey_local_56_sva_1, RoundKey_local_57_sva_1,
      RoundKey_local_58_sva_1, RoundKey_local_59_sva_1, RoundKey_local_60_sva_1,
      RoundKey_local_61_sva_1, RoundKey_local_62_sva_1, RoundKey_local_63_sva_1,
      RoundKey_local_64_sva_1, RoundKey_local_65_sva_1, RoundKey_local_66_sva_1,
      RoundKey_local_67_sva_1, RoundKey_local_68_sva_1, RoundKey_local_69_sva_1,
      RoundKey_local_70_sva_1, RoundKey_local_71_sva_1, RoundKey_local_72_sva_1,
      RoundKey_local_73_sva_1, RoundKey_local_74_sva_1, RoundKey_local_75_sva_1,
      RoundKey_local_76_sva_1, RoundKey_local_77_sva_1, RoundKey_local_78_sva_1,
      RoundKey_local_79_sva_1, RoundKey_local_80_sva_1, RoundKey_local_81_sva_1,
      RoundKey_local_82_sva_1, RoundKey_local_83_sva_1, RoundKey_local_84_sva_1,
      RoundKey_local_85_sva_1, RoundKey_local_86_sva_1, RoundKey_local_87_sva_1,
      RoundKey_local_88_sva_1, RoundKey_local_89_sva_1, RoundKey_local_90_sva_1,
      RoundKey_local_91_sva_1, RoundKey_local_92_sva_1, RoundKey_local_93_sva_1,
      RoundKey_local_94_sva_1, RoundKey_local_95_sva_1, RoundKey_local_96_sva_1,
      RoundKey_local_97_sva_1, RoundKey_local_98_sva_1, RoundKey_local_99_sva_1,
      RoundKey_local_100_sva_1, RoundKey_local_101_sva_1, RoundKey_local_102_sva_1,
      RoundKey_local_103_sva_1, RoundKey_local_104_sva_1, RoundKey_local_105_sva_1,
      RoundKey_local_106_sva_1, RoundKey_local_107_sva_1, RoundKey_local_108_sva_1,
      RoundKey_local_109_sva_1, RoundKey_local_110_sva_1, RoundKey_local_111_sva_1,
      RoundKey_local_112_sva_1, RoundKey_local_113_sva_1, RoundKey_local_114_sva_1,
      RoundKey_local_115_sva_1, RoundKey_local_116_sva_1, RoundKey_local_117_sva_1,
      RoundKey_local_118_sva_1, RoundKey_local_119_sva_1, RoundKey_local_120_sva_1,
      RoundKey_local_121_sva_1, RoundKey_local_122_sva_1, RoundKey_local_123_sva_1,
      RoundKey_local_124_sva_1, RoundKey_local_125_sva_1, RoundKey_local_126_sva_1,
      RoundKey_local_127_sva_1, RoundKey_local_128_sva_1, RoundKey_local_129_sva_1,
      RoundKey_local_130_sva_1, RoundKey_local_131_sva_1, RoundKey_local_132_sva_1,
      RoundKey_local_133_sva_1, RoundKey_local_134_sva_1, RoundKey_local_135_sva_1,
      RoundKey_local_136_sva_1, RoundKey_local_137_sva_1, RoundKey_local_138_sva_1,
      RoundKey_local_139_sva_1, RoundKey_local_140_sva_1, RoundKey_local_141_sva_1,
      RoundKey_local_142_sva_1, RoundKey_local_143_sva_1, RoundKey_local_144_sva_1,
      RoundKey_local_145_sva_1, RoundKey_local_146_sva_1, RoundKey_local_147_sva_1,
      RoundKey_local_148_sva_1, RoundKey_local_149_sva_1, RoundKey_local_150_sva_1,
      RoundKey_local_151_sva_1, RoundKey_local_152_sva_1, RoundKey_local_153_sva_1,
      RoundKey_local_154_sva_1, RoundKey_local_155_sva_1, RoundKey_local_156_sva_1,
      RoundKey_local_157_sva_1, RoundKey_local_158_sva_1, RoundKey_local_159_sva_1,
      RoundKey_local_160_sva_1, RoundKey_local_161_sva_1, RoundKey_local_162_sva_1,
      RoundKey_local_163_sva_1, RoundKey_local_164_sva_1, RoundKey_local_165_sva_1,
      RoundKey_local_166_sva_1, RoundKey_local_167_sva_1, RoundKey_local_168_sva_1,
      RoundKey_local_169_sva_1, RoundKey_local_170_sva_1, RoundKey_local_171_sva_1,
      RoundKey_local_172_sva_1, RoundKey_local_173_sva_1, RoundKey_local_174_sva_1,
      for_slc_i_1_8_7_0_ctmp_sva, {round_3_0_sva , i_2_0_sva_1_0 , j_2_0_sva_1_0});
  assign for_1_for_for_1_for_xor_1_cmx_sva_1 = for_1_for_mux_16_nl ^ for_1_for_mux_17_nl;
  assign nl_for_acc_nl = conv_u2u_4_5(z_out[7:4]) + 5'b10101;
  assign for_acc_nl = nl_for_acc_nl[4:0];
  assign for_acc_itm_4 = readslicef_5_1_4(for_acc_nl);
  assign or_dcpl_1 = (z_out[3:2]!=2'b00);
  assign or_dcpl_2 = (z_out[1:0]!=2'b00);
  assign or_dcpl_3 = or_dcpl_2 | or_dcpl_1;
  assign or_dcpl_4 = (z_out[5:4]!=2'b00);
  assign or_dcpl_5 = (~ for_acc_itm_4) | (z_out[6]);
  assign or_dcpl_6 = or_dcpl_5 | (z_out[7]);
  assign or_dcpl_7 = or_dcpl_6 | or_dcpl_4;
  assign or_dcpl_9 = (z_out[1:0]!=2'b01);
  assign or_dcpl_10 = or_dcpl_9 | or_dcpl_1;
  assign or_dcpl_12 = (z_out[1:0]!=2'b10);
  assign or_dcpl_13 = or_dcpl_12 | or_dcpl_1;
  assign or_dcpl_15 = ~((z_out[1:0]==2'b11));
  assign or_dcpl_16 = or_dcpl_15 | or_dcpl_1;
  assign or_dcpl_18 = (z_out[3:2]!=2'b01);
  assign or_dcpl_19 = or_dcpl_2 | or_dcpl_18;
  assign or_dcpl_21 = or_dcpl_9 | or_dcpl_18;
  assign or_dcpl_23 = or_dcpl_12 | or_dcpl_18;
  assign or_dcpl_25 = or_dcpl_15 | or_dcpl_18;
  assign or_dcpl_27 = (z_out[3:2]!=2'b10);
  assign or_dcpl_28 = or_dcpl_2 | or_dcpl_27;
  assign or_dcpl_30 = or_dcpl_9 | or_dcpl_27;
  assign or_dcpl_32 = or_dcpl_12 | or_dcpl_27;
  assign or_dcpl_34 = or_dcpl_15 | or_dcpl_27;
  assign or_dcpl_36 = ~((z_out[3:2]==2'b11));
  assign or_dcpl_37 = or_dcpl_2 | or_dcpl_36;
  assign or_dcpl_39 = or_dcpl_9 | or_dcpl_36;
  assign or_dcpl_41 = or_dcpl_12 | or_dcpl_36;
  assign or_dcpl_43 = or_dcpl_15 | or_dcpl_36;
  assign or_dcpl_45 = (z_out[5:4]!=2'b01);
  assign or_dcpl_46 = or_dcpl_6 | or_dcpl_45;
  assign or_dcpl_63 = (z_out[5:4]!=2'b10);
  assign or_dcpl_64 = or_dcpl_6 | or_dcpl_63;
  assign or_dcpl_81 = ~((z_out[5:4]==2'b11));
  assign or_dcpl_82 = or_dcpl_6 | or_dcpl_81;
  assign or_dcpl_100 = (~ for_acc_itm_4) | (z_out[7:6]!=2'b01);
  assign or_dcpl_101 = or_dcpl_100 | or_dcpl_4;
  assign or_dcpl_118 = or_dcpl_100 | or_dcpl_45;
  assign or_dcpl_135 = or_dcpl_100 | or_dcpl_63;
  assign or_dcpl_152 = or_dcpl_100 | or_dcpl_81;
  assign or_dcpl_169 = or_dcpl_5 | (~ (z_out[7]));
  assign or_dcpl_170 = or_dcpl_169 | or_dcpl_4;
  assign or_dcpl_187 = or_dcpl_169 | or_dcpl_45;
  assign or_dcpl_204 = or_dcpl_169 | or_dcpl_63;
  assign or_dcpl_224 = (for_slc_i_1_8_7_0_ctmp_sva[1:0]!=2'b00);
  assign or_dcpl_225 = (for_slc_i_1_8_7_0_ctmp_sva[3:2]!=2'b00);
  assign or_dcpl_226 = or_dcpl_225 | or_dcpl_224;
  assign or_dcpl_227 = (for_slc_i_1_8_7_0_ctmp_sva[5:4]!=2'b00);
  assign or_dcpl_228 = (for_slc_i_1_8_7_0_ctmp_sva[7:6]!=2'b00);
  assign or_dcpl_229 = or_dcpl_228 | or_dcpl_227;
  assign or_dcpl_231 = (for_slc_i_1_8_7_0_ctmp_sva[1:0]!=2'b01);
  assign or_dcpl_232 = or_dcpl_225 | or_dcpl_231;
  assign or_dcpl_234 = (for_slc_i_1_8_7_0_ctmp_sva[1:0]!=2'b10);
  assign or_dcpl_235 = or_dcpl_225 | or_dcpl_234;
  assign or_dcpl_237 = ~((for_slc_i_1_8_7_0_ctmp_sva[1:0]==2'b11));
  assign or_dcpl_238 = or_dcpl_225 | or_dcpl_237;
  assign or_dcpl_240 = (for_slc_i_1_8_7_0_ctmp_sva[3:2]!=2'b01);
  assign or_dcpl_241 = or_dcpl_240 | or_dcpl_224;
  assign or_dcpl_243 = or_dcpl_240 | or_dcpl_231;
  assign or_dcpl_245 = or_dcpl_240 | or_dcpl_234;
  assign or_dcpl_247 = or_dcpl_240 | or_dcpl_237;
  assign or_dcpl_249 = (for_slc_i_1_8_7_0_ctmp_sva[3:2]!=2'b10);
  assign or_dcpl_250 = or_dcpl_249 | or_dcpl_224;
  assign or_dcpl_252 = or_dcpl_249 | or_dcpl_231;
  assign or_dcpl_254 = or_dcpl_249 | or_dcpl_234;
  assign or_dcpl_256 = or_dcpl_249 | or_dcpl_237;
  assign or_dcpl_258 = ~((for_slc_i_1_8_7_0_ctmp_sva[3:2]==2'b11));
  assign or_dcpl_259 = or_dcpl_258 | or_dcpl_224;
  assign or_dcpl_261 = or_dcpl_258 | or_dcpl_231;
  assign or_dcpl_263 = or_dcpl_258 | or_dcpl_234;
  assign or_dcpl_265 = or_dcpl_258 | or_dcpl_237;
  assign or_dcpl_267 = (for_slc_i_1_8_7_0_ctmp_sva[5:4]!=2'b01);
  assign or_dcpl_268 = or_dcpl_228 | or_dcpl_267;
  assign or_dcpl_285 = (for_slc_i_1_8_7_0_ctmp_sva[5:4]!=2'b10);
  assign or_dcpl_286 = or_dcpl_228 | or_dcpl_285;
  assign or_dcpl_303 = ~((for_slc_i_1_8_7_0_ctmp_sva[5:4]==2'b11));
  assign or_dcpl_304 = or_dcpl_228 | or_dcpl_303;
  assign or_dcpl_321 = (for_slc_i_1_8_7_0_ctmp_sva[7:6]!=2'b01);
  assign or_dcpl_322 = or_dcpl_321 | or_dcpl_227;
  assign or_dcpl_339 = or_dcpl_321 | or_dcpl_267;
  assign or_dcpl_356 = or_dcpl_321 | or_dcpl_285;
  assign or_dcpl_373 = or_dcpl_321 | or_dcpl_303;
  assign or_dcpl_390 = (for_slc_i_1_8_7_0_ctmp_sva[7:6]!=2'b10);
  assign or_dcpl_391 = or_dcpl_390 | or_dcpl_227;
  assign or_dcpl_408 = or_dcpl_390 | or_dcpl_267;
  assign or_dcpl_425 = or_dcpl_390 | or_dcpl_285;
  assign or_dcpl_441 = (i_2_0_sva_1_0!=2'b00);
  assign or_dcpl_442 = (j_2_0_sva_1_0!=2'b01);
  assign or_dcpl_444 = (j_2_0_sva_1_0!=2'b10);
  assign or_dcpl_446 = ~((j_2_0_sva_1_0==2'b11));
  assign or_dcpl_448 = (i_2_0_sva_1_0!=2'b01);
  assign or_dcpl_449 = (j_2_0_sva_1_0!=2'b00);
  assign or_dcpl_454 = (i_2_0_sva_1_0!=2'b10);
  assign or_dcpl_459 = ~((i_2_0_sva_1_0==2'b11));
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_0_sva_1 <= 8'b00000000;
    end
    else if ( ~(or_dcpl_229 | or_dcpl_226 | (fsm_output[4:2]!=3'b000)) ) begin
      RoundKey_local_0_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_1_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_10) & (~(or_dcpl_229 | or_dcpl_232))
        ) begin
      RoundKey_local_1_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_2_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_13) & (~(or_dcpl_229 | or_dcpl_235))
        ) begin
      RoundKey_local_2_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_3_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_16) & (~(or_dcpl_229 | or_dcpl_238))
        ) begin
      RoundKey_local_3_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_4_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_19) & (~(or_dcpl_229 | or_dcpl_241))
        ) begin
      RoundKey_local_4_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_5_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_21) & (~(or_dcpl_229 | or_dcpl_243))
        ) begin
      RoundKey_local_5_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_6_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_23) & (~(or_dcpl_229 | or_dcpl_245))
        ) begin
      RoundKey_local_6_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_7_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_25) & (~(or_dcpl_229 | or_dcpl_247))
        ) begin
      RoundKey_local_7_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_8_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_28) & (~(or_dcpl_229 | or_dcpl_250))
        ) begin
      RoundKey_local_8_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_9_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_30) & (~(or_dcpl_229 | or_dcpl_252))
        ) begin
      RoundKey_local_9_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_10_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_32) & (~(or_dcpl_229 | or_dcpl_254))
        ) begin
      RoundKey_local_10_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_11_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_34) & (~(or_dcpl_229 | or_dcpl_256))
        ) begin
      RoundKey_local_11_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_12_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_37) & (~(or_dcpl_229 | or_dcpl_259))
        ) begin
      RoundKey_local_12_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_13_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_39) & (~(or_dcpl_229 | or_dcpl_261))
        ) begin
      RoundKey_local_13_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_14_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_41) & (~(or_dcpl_229 | or_dcpl_263))
        ) begin
      RoundKey_local_14_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_15_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_7 | or_dcpl_43) & (~(or_dcpl_229 | or_dcpl_265))
        ) begin
      RoundKey_local_15_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_16_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_3) & (~(or_dcpl_268 | or_dcpl_226))
        ) begin
      RoundKey_local_16_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_17_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_10) & (~(or_dcpl_268 | or_dcpl_232))
        ) begin
      RoundKey_local_17_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_18_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_13) & (~(or_dcpl_268 | or_dcpl_235))
        ) begin
      RoundKey_local_18_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_19_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_16) & (~(or_dcpl_268 | or_dcpl_238))
        ) begin
      RoundKey_local_19_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_20_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_19) & (~(or_dcpl_268 | or_dcpl_241))
        ) begin
      RoundKey_local_20_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_21_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_21) & (~(or_dcpl_268 | or_dcpl_243))
        ) begin
      RoundKey_local_21_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_22_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_23) & (~(or_dcpl_268 | or_dcpl_245))
        ) begin
      RoundKey_local_22_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_23_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_25) & (~(or_dcpl_268 | or_dcpl_247))
        ) begin
      RoundKey_local_23_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_24_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_28) & (~(or_dcpl_268 | or_dcpl_250))
        ) begin
      RoundKey_local_24_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_25_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_30) & (~(or_dcpl_268 | or_dcpl_252))
        ) begin
      RoundKey_local_25_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_26_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_32) & (~(or_dcpl_268 | or_dcpl_254))
        ) begin
      RoundKey_local_26_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_27_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_34) & (~(or_dcpl_268 | or_dcpl_256))
        ) begin
      RoundKey_local_27_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_28_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_37) & (~(or_dcpl_268 | or_dcpl_259))
        ) begin
      RoundKey_local_28_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_29_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_39) & (~(or_dcpl_268 | or_dcpl_261))
        ) begin
      RoundKey_local_29_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_30_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_41) & (~(or_dcpl_268 | or_dcpl_263))
        ) begin
      RoundKey_local_30_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_31_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_46 | or_dcpl_43) & (~(or_dcpl_268 | or_dcpl_265))
        ) begin
      RoundKey_local_31_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_32_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_3) & (~(or_dcpl_286 | or_dcpl_226))
        ) begin
      RoundKey_local_32_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_33_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_10) & (~(or_dcpl_286 | or_dcpl_232))
        ) begin
      RoundKey_local_33_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_34_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_13) & (~(or_dcpl_286 | or_dcpl_235))
        ) begin
      RoundKey_local_34_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_35_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_16) & (~(or_dcpl_286 | or_dcpl_238))
        ) begin
      RoundKey_local_35_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_36_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_19) & (~(or_dcpl_286 | or_dcpl_241))
        ) begin
      RoundKey_local_36_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_37_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_21) & (~(or_dcpl_286 | or_dcpl_243))
        ) begin
      RoundKey_local_37_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_38_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_23) & (~(or_dcpl_286 | or_dcpl_245))
        ) begin
      RoundKey_local_38_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_39_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_25) & (~(or_dcpl_286 | or_dcpl_247))
        ) begin
      RoundKey_local_39_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_40_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_28) & (~(or_dcpl_286 | or_dcpl_250))
        ) begin
      RoundKey_local_40_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_41_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_30) & (~(or_dcpl_286 | or_dcpl_252))
        ) begin
      RoundKey_local_41_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_42_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_32) & (~(or_dcpl_286 | or_dcpl_254))
        ) begin
      RoundKey_local_42_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_43_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_34) & (~(or_dcpl_286 | or_dcpl_256))
        ) begin
      RoundKey_local_43_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_44_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_37) & (~(or_dcpl_286 | or_dcpl_259))
        ) begin
      RoundKey_local_44_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_45_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_39) & (~(or_dcpl_286 | or_dcpl_261))
        ) begin
      RoundKey_local_45_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_46_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_41) & (~(or_dcpl_286 | or_dcpl_263))
        ) begin
      RoundKey_local_46_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_47_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_64 | or_dcpl_43) & (~(or_dcpl_286 | or_dcpl_265))
        ) begin
      RoundKey_local_47_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_48_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_3) & (~(or_dcpl_304 | or_dcpl_226))
        ) begin
      RoundKey_local_48_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_49_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_10) & (~(or_dcpl_304 | or_dcpl_232))
        ) begin
      RoundKey_local_49_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_50_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_13) & (~(or_dcpl_304 | or_dcpl_235))
        ) begin
      RoundKey_local_50_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_51_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_16) & (~(or_dcpl_304 | or_dcpl_238))
        ) begin
      RoundKey_local_51_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_52_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_19) & (~(or_dcpl_304 | or_dcpl_241))
        ) begin
      RoundKey_local_52_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_53_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_21) & (~(or_dcpl_304 | or_dcpl_243))
        ) begin
      RoundKey_local_53_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_54_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_23) & (~(or_dcpl_304 | or_dcpl_245))
        ) begin
      RoundKey_local_54_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_55_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_25) & (~(or_dcpl_304 | or_dcpl_247))
        ) begin
      RoundKey_local_55_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_56_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_28) & (~(or_dcpl_304 | or_dcpl_250))
        ) begin
      RoundKey_local_56_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_57_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_30) & (~(or_dcpl_304 | or_dcpl_252))
        ) begin
      RoundKey_local_57_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_58_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_32) & (~(or_dcpl_304 | or_dcpl_254))
        ) begin
      RoundKey_local_58_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_59_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_34) & (~(or_dcpl_304 | or_dcpl_256))
        ) begin
      RoundKey_local_59_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_60_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_37) & (~(or_dcpl_304 | or_dcpl_259))
        ) begin
      RoundKey_local_60_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_61_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_39) & (~(or_dcpl_304 | or_dcpl_261))
        ) begin
      RoundKey_local_61_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_62_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_41) & (~(or_dcpl_304 | or_dcpl_263))
        ) begin
      RoundKey_local_62_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_63_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_82 | or_dcpl_43) & (~(or_dcpl_304 | or_dcpl_265))
        ) begin
      RoundKey_local_63_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_64_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_3) & (~(or_dcpl_322 | or_dcpl_226))
        ) begin
      RoundKey_local_64_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_65_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_10) & (~(or_dcpl_322 | or_dcpl_232))
        ) begin
      RoundKey_local_65_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_66_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_13) & (~(or_dcpl_322 | or_dcpl_235))
        ) begin
      RoundKey_local_66_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_67_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_16) & (~(or_dcpl_322 | or_dcpl_238))
        ) begin
      RoundKey_local_67_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_68_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_19) & (~(or_dcpl_322 | or_dcpl_241))
        ) begin
      RoundKey_local_68_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_69_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_21) & (~(or_dcpl_322 | or_dcpl_243))
        ) begin
      RoundKey_local_69_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_70_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_23) & (~(or_dcpl_322 | or_dcpl_245))
        ) begin
      RoundKey_local_70_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_71_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_25) & (~(or_dcpl_322 | or_dcpl_247))
        ) begin
      RoundKey_local_71_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_72_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_28) & (~(or_dcpl_322 | or_dcpl_250))
        ) begin
      RoundKey_local_72_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_73_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_30) & (~(or_dcpl_322 | or_dcpl_252))
        ) begin
      RoundKey_local_73_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_74_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_32) & (~(or_dcpl_322 | or_dcpl_254))
        ) begin
      RoundKey_local_74_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_75_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_34) & (~(or_dcpl_322 | or_dcpl_256))
        ) begin
      RoundKey_local_75_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_76_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_37) & (~(or_dcpl_322 | or_dcpl_259))
        ) begin
      RoundKey_local_76_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_77_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_39) & (~(or_dcpl_322 | or_dcpl_261))
        ) begin
      RoundKey_local_77_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_78_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_41) & (~(or_dcpl_322 | or_dcpl_263))
        ) begin
      RoundKey_local_78_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_79_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_101 | or_dcpl_43) & (~(or_dcpl_322 | or_dcpl_265))
        ) begin
      RoundKey_local_79_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_80_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_3) & (~(or_dcpl_339 | or_dcpl_226))
        ) begin
      RoundKey_local_80_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_81_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_10) & (~(or_dcpl_339 | or_dcpl_232))
        ) begin
      RoundKey_local_81_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_82_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_13) & (~(or_dcpl_339 | or_dcpl_235))
        ) begin
      RoundKey_local_82_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_83_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_16) & (~(or_dcpl_339 | or_dcpl_238))
        ) begin
      RoundKey_local_83_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_84_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_19) & (~(or_dcpl_339 | or_dcpl_241))
        ) begin
      RoundKey_local_84_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_85_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_21) & (~(or_dcpl_339 | or_dcpl_243))
        ) begin
      RoundKey_local_85_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_86_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_23) & (~(or_dcpl_339 | or_dcpl_245))
        ) begin
      RoundKey_local_86_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_87_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_25) & (~(or_dcpl_339 | or_dcpl_247))
        ) begin
      RoundKey_local_87_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_88_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_28) & (~(or_dcpl_339 | or_dcpl_250))
        ) begin
      RoundKey_local_88_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_89_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_30) & (~(or_dcpl_339 | or_dcpl_252))
        ) begin
      RoundKey_local_89_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_90_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_32) & (~(or_dcpl_339 | or_dcpl_254))
        ) begin
      RoundKey_local_90_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_91_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_34) & (~(or_dcpl_339 | or_dcpl_256))
        ) begin
      RoundKey_local_91_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_92_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_37) & (~(or_dcpl_339 | or_dcpl_259))
        ) begin
      RoundKey_local_92_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_93_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_39) & (~(or_dcpl_339 | or_dcpl_261))
        ) begin
      RoundKey_local_93_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_94_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_41) & (~(or_dcpl_339 | or_dcpl_263))
        ) begin
      RoundKey_local_94_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_95_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_118 | or_dcpl_43) & (~(or_dcpl_339 | or_dcpl_265))
        ) begin
      RoundKey_local_95_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_96_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_3) & (~(or_dcpl_356 | or_dcpl_226))
        ) begin
      RoundKey_local_96_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_97_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_10) & (~(or_dcpl_356 | or_dcpl_232))
        ) begin
      RoundKey_local_97_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_98_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_13) & (~(or_dcpl_356 | or_dcpl_235))
        ) begin
      RoundKey_local_98_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_99_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_16) & (~(or_dcpl_356 | or_dcpl_238))
        ) begin
      RoundKey_local_99_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_100_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_19) & (~(or_dcpl_356 | or_dcpl_241))
        ) begin
      RoundKey_local_100_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_101_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_21) & (~(or_dcpl_356 | or_dcpl_243))
        ) begin
      RoundKey_local_101_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_102_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_23) & (~(or_dcpl_356 | or_dcpl_245))
        ) begin
      RoundKey_local_102_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_103_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_25) & (~(or_dcpl_356 | or_dcpl_247))
        ) begin
      RoundKey_local_103_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_104_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_28) & (~(or_dcpl_356 | or_dcpl_250))
        ) begin
      RoundKey_local_104_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_105_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_30) & (~(or_dcpl_356 | or_dcpl_252))
        ) begin
      RoundKey_local_105_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_106_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_32) & (~(or_dcpl_356 | or_dcpl_254))
        ) begin
      RoundKey_local_106_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_107_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_34) & (~(or_dcpl_356 | or_dcpl_256))
        ) begin
      RoundKey_local_107_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_108_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_37) & (~(or_dcpl_356 | or_dcpl_259))
        ) begin
      RoundKey_local_108_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_109_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_39) & (~(or_dcpl_356 | or_dcpl_261))
        ) begin
      RoundKey_local_109_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_110_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_41) & (~(or_dcpl_356 | or_dcpl_263))
        ) begin
      RoundKey_local_110_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_111_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_135 | or_dcpl_43) & (~(or_dcpl_356 | or_dcpl_265))
        ) begin
      RoundKey_local_111_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_112_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_3) & (~(or_dcpl_373 | or_dcpl_226))
        ) begin
      RoundKey_local_112_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_113_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_10) & (~(or_dcpl_373 | or_dcpl_232))
        ) begin
      RoundKey_local_113_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_114_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_13) & (~(or_dcpl_373 | or_dcpl_235))
        ) begin
      RoundKey_local_114_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_115_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_16) & (~(or_dcpl_373 | or_dcpl_238))
        ) begin
      RoundKey_local_115_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_116_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_19) & (~(or_dcpl_373 | or_dcpl_241))
        ) begin
      RoundKey_local_116_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_117_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_21) & (~(or_dcpl_373 | or_dcpl_243))
        ) begin
      RoundKey_local_117_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_118_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_23) & (~(or_dcpl_373 | or_dcpl_245))
        ) begin
      RoundKey_local_118_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_119_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_25) & (~(or_dcpl_373 | or_dcpl_247))
        ) begin
      RoundKey_local_119_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_120_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_28) & (~(or_dcpl_373 | or_dcpl_250))
        ) begin
      RoundKey_local_120_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_121_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_30) & (~(or_dcpl_373 | or_dcpl_252))
        ) begin
      RoundKey_local_121_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_122_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_32) & (~(or_dcpl_373 | or_dcpl_254))
        ) begin
      RoundKey_local_122_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_123_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_34) & (~(or_dcpl_373 | or_dcpl_256))
        ) begin
      RoundKey_local_123_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_124_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_37) & (~(or_dcpl_373 | or_dcpl_259))
        ) begin
      RoundKey_local_124_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_125_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_39) & (~(or_dcpl_373 | or_dcpl_261))
        ) begin
      RoundKey_local_125_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_126_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_41) & (~(or_dcpl_373 | or_dcpl_263))
        ) begin
      RoundKey_local_126_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_127_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_152 | or_dcpl_43) & (~(or_dcpl_373 | or_dcpl_265))
        ) begin
      RoundKey_local_127_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_128_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_3) & (~(or_dcpl_391 | or_dcpl_226))
        ) begin
      RoundKey_local_128_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_129_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_10) & (~(or_dcpl_391 | or_dcpl_232))
        ) begin
      RoundKey_local_129_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_130_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_13) & (~(or_dcpl_391 | or_dcpl_235))
        ) begin
      RoundKey_local_130_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_131_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_16) & (~(or_dcpl_391 | or_dcpl_238))
        ) begin
      RoundKey_local_131_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_132_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_19) & (~(or_dcpl_391 | or_dcpl_241))
        ) begin
      RoundKey_local_132_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_133_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_21) & (~(or_dcpl_391 | or_dcpl_243))
        ) begin
      RoundKey_local_133_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_134_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_23) & (~(or_dcpl_391 | or_dcpl_245))
        ) begin
      RoundKey_local_134_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_135_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_25) & (~(or_dcpl_391 | or_dcpl_247))
        ) begin
      RoundKey_local_135_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_136_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_28) & (~(or_dcpl_391 | or_dcpl_250))
        ) begin
      RoundKey_local_136_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_137_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_30) & (~(or_dcpl_391 | or_dcpl_252))
        ) begin
      RoundKey_local_137_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_138_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_32) & (~(or_dcpl_391 | or_dcpl_254))
        ) begin
      RoundKey_local_138_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_139_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_34) & (~(or_dcpl_391 | or_dcpl_256))
        ) begin
      RoundKey_local_139_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_140_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_37) & (~(or_dcpl_391 | or_dcpl_259))
        ) begin
      RoundKey_local_140_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_141_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_39) & (~(or_dcpl_391 | or_dcpl_261))
        ) begin
      RoundKey_local_141_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_142_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_41) & (~(or_dcpl_391 | or_dcpl_263))
        ) begin
      RoundKey_local_142_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_143_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_170 | or_dcpl_43) & (~(or_dcpl_391 | or_dcpl_265))
        ) begin
      RoundKey_local_143_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_144_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_3) & (~(or_dcpl_408 | or_dcpl_226))
        ) begin
      RoundKey_local_144_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_145_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_10) & (~(or_dcpl_408 | or_dcpl_232))
        ) begin
      RoundKey_local_145_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_146_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_13) & (~(or_dcpl_408 | or_dcpl_235))
        ) begin
      RoundKey_local_146_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_147_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_16) & (~(or_dcpl_408 | or_dcpl_238))
        ) begin
      RoundKey_local_147_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_148_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_19) & (~(or_dcpl_408 | or_dcpl_241))
        ) begin
      RoundKey_local_148_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_149_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_21) & (~(or_dcpl_408 | or_dcpl_243))
        ) begin
      RoundKey_local_149_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_150_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_23) & (~(or_dcpl_408 | or_dcpl_245))
        ) begin
      RoundKey_local_150_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_151_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_25) & (~(or_dcpl_408 | or_dcpl_247))
        ) begin
      RoundKey_local_151_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_152_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_28) & (~(or_dcpl_408 | or_dcpl_250))
        ) begin
      RoundKey_local_152_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_153_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_30) & (~(or_dcpl_408 | or_dcpl_252))
        ) begin
      RoundKey_local_153_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_154_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_32) & (~(or_dcpl_408 | or_dcpl_254))
        ) begin
      RoundKey_local_154_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_155_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_34) & (~(or_dcpl_408 | or_dcpl_256))
        ) begin
      RoundKey_local_155_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_156_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_37) & (~(or_dcpl_408 | or_dcpl_259))
        ) begin
      RoundKey_local_156_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_157_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_39) & (~(or_dcpl_408 | or_dcpl_261))
        ) begin
      RoundKey_local_157_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_158_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_41) & (~(or_dcpl_408 | or_dcpl_263))
        ) begin
      RoundKey_local_158_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_159_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_187 | or_dcpl_43) & (~(or_dcpl_408 | or_dcpl_265))
        ) begin
      RoundKey_local_159_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_160_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_3) & (~(or_dcpl_425 | or_dcpl_226))
        ) begin
      RoundKey_local_160_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_161_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_10) & (~(or_dcpl_425 | or_dcpl_232))
        ) begin
      RoundKey_local_161_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_162_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_13) & (~(or_dcpl_425 | or_dcpl_235))
        ) begin
      RoundKey_local_162_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_163_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_16) & (~(or_dcpl_425 | or_dcpl_238))
        ) begin
      RoundKey_local_163_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_164_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_19) & (~(or_dcpl_425 | or_dcpl_241))
        ) begin
      RoundKey_local_164_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_165_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_21) & (~(or_dcpl_425 | or_dcpl_243))
        ) begin
      RoundKey_local_165_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_166_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_23) & (~(or_dcpl_425 | or_dcpl_245))
        ) begin
      RoundKey_local_166_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_167_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_25) & (~(or_dcpl_425 | or_dcpl_247))
        ) begin
      RoundKey_local_167_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_168_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_28) & (~(or_dcpl_425 | or_dcpl_250))
        ) begin
      RoundKey_local_168_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_169_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_30) & (~(or_dcpl_425 | or_dcpl_252))
        ) begin
      RoundKey_local_169_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_170_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_32) & (~(or_dcpl_425 | or_dcpl_254))
        ) begin
      RoundKey_local_170_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_171_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_34) & (~(or_dcpl_425 | or_dcpl_256))
        ) begin
      RoundKey_local_171_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_172_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_37) & (~(or_dcpl_425 | or_dcpl_259))
        ) begin
      RoundKey_local_172_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_173_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_39) & (~(or_dcpl_425 | or_dcpl_261))
        ) begin
      RoundKey_local_173_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      RoundKey_local_174_sva_1 <= 8'b00000000;
    end
    else if ( (fsm_output[1]) & (or_dcpl_204 | or_dcpl_41) & (~(or_dcpl_425 | or_dcpl_263))
        ) begin
      RoundKey_local_174_sva_1 <= for_slc_i_1_8_7_0_ctmp_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      round_3_0_sva <= 4'b0000;
    end
    else if ( ~ nor_rgt ) begin
      round_3_0_sva <= round_rsci_idat[3:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      reg_RoundKey_triosy_obj_ld_cse <= 1'b0;
    end
    else begin
      reg_RoundKey_triosy_obj_ld_cse <= (z_out[2]) & (fsm_output[4]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      for_slc_i_1_8_7_0_ctmp_sva <= 8'b00000000;
    end
    else if ( (fsm_output[5]) | (fsm_output[0]) | (fsm_output[1]) ) begin
      for_slc_i_1_8_7_0_ctmp_sva <= MUX_v_8_2_2(8'b00000000, for_for_mux_nl, nor_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      i_2_0_sva_1_0 <= 2'b00;
    end
    else if ( (fsm_output[4]) | (fsm_output[1]) ) begin
      i_2_0_sva_1_0 <= MUX_v_2_2_2(2'b00, (z_out[1:0]), (fsm_output[4]));
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      j_2_0_sva_1_0 <= 2'b00;
    end
    else if ( (fsm_output[4]) | (fsm_output[1]) | (fsm_output[3]) ) begin
      j_2_0_sva_1_0 <= MUX_v_2_2_2(2'b00, (z_out[1:0]), (fsm_output[3]));
    end
  end
  assign and_372_nl = for_acc_itm_4 & (fsm_output[1]);
  assign for_for_mux_nl = MUX_v_8_2_2(for_slc_i_1_8_7_0_ctmp_sva_mx0w1, z_out, and_372_nl);
  assign for_nor_2_nl = ~((fsm_output[4:3]!=2'b00));
  assign for_for_and_1_nl = MUX_v_6_2_2(6'b000000, (for_slc_i_1_8_7_0_ctmp_sva[7:2]),
      for_nor_2_nl);
  assign for_mux1h_3_nl = MUX1HOT_v_2_3_2((for_slc_i_1_8_7_0_ctmp_sva[1:0]), j_2_0_sva_1_0,
      i_2_0_sva_1_0, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_z_out = ({for_for_and_1_nl , for_mux1h_3_nl}) + 8'b00000001;
  assign z_out = nl_z_out[7:0];

  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_16_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [3:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_8_16_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_176_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [7:0] input_16;
    input [7:0] input_17;
    input [7:0] input_18;
    input [7:0] input_19;
    input [7:0] input_20;
    input [7:0] input_21;
    input [7:0] input_22;
    input [7:0] input_23;
    input [7:0] input_24;
    input [7:0] input_25;
    input [7:0] input_26;
    input [7:0] input_27;
    input [7:0] input_28;
    input [7:0] input_29;
    input [7:0] input_30;
    input [7:0] input_31;
    input [7:0] input_32;
    input [7:0] input_33;
    input [7:0] input_34;
    input [7:0] input_35;
    input [7:0] input_36;
    input [7:0] input_37;
    input [7:0] input_38;
    input [7:0] input_39;
    input [7:0] input_40;
    input [7:0] input_41;
    input [7:0] input_42;
    input [7:0] input_43;
    input [7:0] input_44;
    input [7:0] input_45;
    input [7:0] input_46;
    input [7:0] input_47;
    input [7:0] input_48;
    input [7:0] input_49;
    input [7:0] input_50;
    input [7:0] input_51;
    input [7:0] input_52;
    input [7:0] input_53;
    input [7:0] input_54;
    input [7:0] input_55;
    input [7:0] input_56;
    input [7:0] input_57;
    input [7:0] input_58;
    input [7:0] input_59;
    input [7:0] input_60;
    input [7:0] input_61;
    input [7:0] input_62;
    input [7:0] input_63;
    input [7:0] input_64;
    input [7:0] input_65;
    input [7:0] input_66;
    input [7:0] input_67;
    input [7:0] input_68;
    input [7:0] input_69;
    input [7:0] input_70;
    input [7:0] input_71;
    input [7:0] input_72;
    input [7:0] input_73;
    input [7:0] input_74;
    input [7:0] input_75;
    input [7:0] input_76;
    input [7:0] input_77;
    input [7:0] input_78;
    input [7:0] input_79;
    input [7:0] input_80;
    input [7:0] input_81;
    input [7:0] input_82;
    input [7:0] input_83;
    input [7:0] input_84;
    input [7:0] input_85;
    input [7:0] input_86;
    input [7:0] input_87;
    input [7:0] input_88;
    input [7:0] input_89;
    input [7:0] input_90;
    input [7:0] input_91;
    input [7:0] input_92;
    input [7:0] input_93;
    input [7:0] input_94;
    input [7:0] input_95;
    input [7:0] input_96;
    input [7:0] input_97;
    input [7:0] input_98;
    input [7:0] input_99;
    input [7:0] input_100;
    input [7:0] input_101;
    input [7:0] input_102;
    input [7:0] input_103;
    input [7:0] input_104;
    input [7:0] input_105;
    input [7:0] input_106;
    input [7:0] input_107;
    input [7:0] input_108;
    input [7:0] input_109;
    input [7:0] input_110;
    input [7:0] input_111;
    input [7:0] input_112;
    input [7:0] input_113;
    input [7:0] input_114;
    input [7:0] input_115;
    input [7:0] input_116;
    input [7:0] input_117;
    input [7:0] input_118;
    input [7:0] input_119;
    input [7:0] input_120;
    input [7:0] input_121;
    input [7:0] input_122;
    input [7:0] input_123;
    input [7:0] input_124;
    input [7:0] input_125;
    input [7:0] input_126;
    input [7:0] input_127;
    input [7:0] input_128;
    input [7:0] input_129;
    input [7:0] input_130;
    input [7:0] input_131;
    input [7:0] input_132;
    input [7:0] input_133;
    input [7:0] input_134;
    input [7:0] input_135;
    input [7:0] input_136;
    input [7:0] input_137;
    input [7:0] input_138;
    input [7:0] input_139;
    input [7:0] input_140;
    input [7:0] input_141;
    input [7:0] input_142;
    input [7:0] input_143;
    input [7:0] input_144;
    input [7:0] input_145;
    input [7:0] input_146;
    input [7:0] input_147;
    input [7:0] input_148;
    input [7:0] input_149;
    input [7:0] input_150;
    input [7:0] input_151;
    input [7:0] input_152;
    input [7:0] input_153;
    input [7:0] input_154;
    input [7:0] input_155;
    input [7:0] input_156;
    input [7:0] input_157;
    input [7:0] input_158;
    input [7:0] input_159;
    input [7:0] input_160;
    input [7:0] input_161;
    input [7:0] input_162;
    input [7:0] input_163;
    input [7:0] input_164;
    input [7:0] input_165;
    input [7:0] input_166;
    input [7:0] input_167;
    input [7:0] input_168;
    input [7:0] input_169;
    input [7:0] input_170;
    input [7:0] input_171;
    input [7:0] input_172;
    input [7:0] input_173;
    input [7:0] input_174;
    input [7:0] input_175;
    input [7:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      8'b00000000 : begin
        result = input_0;
      end
      8'b00000001 : begin
        result = input_1;
      end
      8'b00000010 : begin
        result = input_2;
      end
      8'b00000011 : begin
        result = input_3;
      end
      8'b00000100 : begin
        result = input_4;
      end
      8'b00000101 : begin
        result = input_5;
      end
      8'b00000110 : begin
        result = input_6;
      end
      8'b00000111 : begin
        result = input_7;
      end
      8'b00001000 : begin
        result = input_8;
      end
      8'b00001001 : begin
        result = input_9;
      end
      8'b00001010 : begin
        result = input_10;
      end
      8'b00001011 : begin
        result = input_11;
      end
      8'b00001100 : begin
        result = input_12;
      end
      8'b00001101 : begin
        result = input_13;
      end
      8'b00001110 : begin
        result = input_14;
      end
      8'b00001111 : begin
        result = input_15;
      end
      8'b00010000 : begin
        result = input_16;
      end
      8'b00010001 : begin
        result = input_17;
      end
      8'b00010010 : begin
        result = input_18;
      end
      8'b00010011 : begin
        result = input_19;
      end
      8'b00010100 : begin
        result = input_20;
      end
      8'b00010101 : begin
        result = input_21;
      end
      8'b00010110 : begin
        result = input_22;
      end
      8'b00010111 : begin
        result = input_23;
      end
      8'b00011000 : begin
        result = input_24;
      end
      8'b00011001 : begin
        result = input_25;
      end
      8'b00011010 : begin
        result = input_26;
      end
      8'b00011011 : begin
        result = input_27;
      end
      8'b00011100 : begin
        result = input_28;
      end
      8'b00011101 : begin
        result = input_29;
      end
      8'b00011110 : begin
        result = input_30;
      end
      8'b00011111 : begin
        result = input_31;
      end
      8'b00100000 : begin
        result = input_32;
      end
      8'b00100001 : begin
        result = input_33;
      end
      8'b00100010 : begin
        result = input_34;
      end
      8'b00100011 : begin
        result = input_35;
      end
      8'b00100100 : begin
        result = input_36;
      end
      8'b00100101 : begin
        result = input_37;
      end
      8'b00100110 : begin
        result = input_38;
      end
      8'b00100111 : begin
        result = input_39;
      end
      8'b00101000 : begin
        result = input_40;
      end
      8'b00101001 : begin
        result = input_41;
      end
      8'b00101010 : begin
        result = input_42;
      end
      8'b00101011 : begin
        result = input_43;
      end
      8'b00101100 : begin
        result = input_44;
      end
      8'b00101101 : begin
        result = input_45;
      end
      8'b00101110 : begin
        result = input_46;
      end
      8'b00101111 : begin
        result = input_47;
      end
      8'b00110000 : begin
        result = input_48;
      end
      8'b00110001 : begin
        result = input_49;
      end
      8'b00110010 : begin
        result = input_50;
      end
      8'b00110011 : begin
        result = input_51;
      end
      8'b00110100 : begin
        result = input_52;
      end
      8'b00110101 : begin
        result = input_53;
      end
      8'b00110110 : begin
        result = input_54;
      end
      8'b00110111 : begin
        result = input_55;
      end
      8'b00111000 : begin
        result = input_56;
      end
      8'b00111001 : begin
        result = input_57;
      end
      8'b00111010 : begin
        result = input_58;
      end
      8'b00111011 : begin
        result = input_59;
      end
      8'b00111100 : begin
        result = input_60;
      end
      8'b00111101 : begin
        result = input_61;
      end
      8'b00111110 : begin
        result = input_62;
      end
      8'b00111111 : begin
        result = input_63;
      end
      8'b01000000 : begin
        result = input_64;
      end
      8'b01000001 : begin
        result = input_65;
      end
      8'b01000010 : begin
        result = input_66;
      end
      8'b01000011 : begin
        result = input_67;
      end
      8'b01000100 : begin
        result = input_68;
      end
      8'b01000101 : begin
        result = input_69;
      end
      8'b01000110 : begin
        result = input_70;
      end
      8'b01000111 : begin
        result = input_71;
      end
      8'b01001000 : begin
        result = input_72;
      end
      8'b01001001 : begin
        result = input_73;
      end
      8'b01001010 : begin
        result = input_74;
      end
      8'b01001011 : begin
        result = input_75;
      end
      8'b01001100 : begin
        result = input_76;
      end
      8'b01001101 : begin
        result = input_77;
      end
      8'b01001110 : begin
        result = input_78;
      end
      8'b01001111 : begin
        result = input_79;
      end
      8'b01010000 : begin
        result = input_80;
      end
      8'b01010001 : begin
        result = input_81;
      end
      8'b01010010 : begin
        result = input_82;
      end
      8'b01010011 : begin
        result = input_83;
      end
      8'b01010100 : begin
        result = input_84;
      end
      8'b01010101 : begin
        result = input_85;
      end
      8'b01010110 : begin
        result = input_86;
      end
      8'b01010111 : begin
        result = input_87;
      end
      8'b01011000 : begin
        result = input_88;
      end
      8'b01011001 : begin
        result = input_89;
      end
      8'b01011010 : begin
        result = input_90;
      end
      8'b01011011 : begin
        result = input_91;
      end
      8'b01011100 : begin
        result = input_92;
      end
      8'b01011101 : begin
        result = input_93;
      end
      8'b01011110 : begin
        result = input_94;
      end
      8'b01011111 : begin
        result = input_95;
      end
      8'b01100000 : begin
        result = input_96;
      end
      8'b01100001 : begin
        result = input_97;
      end
      8'b01100010 : begin
        result = input_98;
      end
      8'b01100011 : begin
        result = input_99;
      end
      8'b01100100 : begin
        result = input_100;
      end
      8'b01100101 : begin
        result = input_101;
      end
      8'b01100110 : begin
        result = input_102;
      end
      8'b01100111 : begin
        result = input_103;
      end
      8'b01101000 : begin
        result = input_104;
      end
      8'b01101001 : begin
        result = input_105;
      end
      8'b01101010 : begin
        result = input_106;
      end
      8'b01101011 : begin
        result = input_107;
      end
      8'b01101100 : begin
        result = input_108;
      end
      8'b01101101 : begin
        result = input_109;
      end
      8'b01101110 : begin
        result = input_110;
      end
      8'b01101111 : begin
        result = input_111;
      end
      8'b01110000 : begin
        result = input_112;
      end
      8'b01110001 : begin
        result = input_113;
      end
      8'b01110010 : begin
        result = input_114;
      end
      8'b01110011 : begin
        result = input_115;
      end
      8'b01110100 : begin
        result = input_116;
      end
      8'b01110101 : begin
        result = input_117;
      end
      8'b01110110 : begin
        result = input_118;
      end
      8'b01110111 : begin
        result = input_119;
      end
      8'b01111000 : begin
        result = input_120;
      end
      8'b01111001 : begin
        result = input_121;
      end
      8'b01111010 : begin
        result = input_122;
      end
      8'b01111011 : begin
        result = input_123;
      end
      8'b01111100 : begin
        result = input_124;
      end
      8'b01111101 : begin
        result = input_125;
      end
      8'b01111110 : begin
        result = input_126;
      end
      8'b01111111 : begin
        result = input_127;
      end
      8'b10000000 : begin
        result = input_128;
      end
      8'b10000001 : begin
        result = input_129;
      end
      8'b10000010 : begin
        result = input_130;
      end
      8'b10000011 : begin
        result = input_131;
      end
      8'b10000100 : begin
        result = input_132;
      end
      8'b10000101 : begin
        result = input_133;
      end
      8'b10000110 : begin
        result = input_134;
      end
      8'b10000111 : begin
        result = input_135;
      end
      8'b10001000 : begin
        result = input_136;
      end
      8'b10001001 : begin
        result = input_137;
      end
      8'b10001010 : begin
        result = input_138;
      end
      8'b10001011 : begin
        result = input_139;
      end
      8'b10001100 : begin
        result = input_140;
      end
      8'b10001101 : begin
        result = input_141;
      end
      8'b10001110 : begin
        result = input_142;
      end
      8'b10001111 : begin
        result = input_143;
      end
      8'b10010000 : begin
        result = input_144;
      end
      8'b10010001 : begin
        result = input_145;
      end
      8'b10010010 : begin
        result = input_146;
      end
      8'b10010011 : begin
        result = input_147;
      end
      8'b10010100 : begin
        result = input_148;
      end
      8'b10010101 : begin
        result = input_149;
      end
      8'b10010110 : begin
        result = input_150;
      end
      8'b10010111 : begin
        result = input_151;
      end
      8'b10011000 : begin
        result = input_152;
      end
      8'b10011001 : begin
        result = input_153;
      end
      8'b10011010 : begin
        result = input_154;
      end
      8'b10011011 : begin
        result = input_155;
      end
      8'b10011100 : begin
        result = input_156;
      end
      8'b10011101 : begin
        result = input_157;
      end
      8'b10011110 : begin
        result = input_158;
      end
      8'b10011111 : begin
        result = input_159;
      end
      8'b10100000 : begin
        result = input_160;
      end
      8'b10100001 : begin
        result = input_161;
      end
      8'b10100010 : begin
        result = input_162;
      end
      8'b10100011 : begin
        result = input_163;
      end
      8'b10100100 : begin
        result = input_164;
      end
      8'b10100101 : begin
        result = input_165;
      end
      8'b10100110 : begin
        result = input_166;
      end
      8'b10100111 : begin
        result = input_167;
      end
      8'b10101000 : begin
        result = input_168;
      end
      8'b10101001 : begin
        result = input_169;
      end
      8'b10101010 : begin
        result = input_170;
      end
      8'b10101011 : begin
        result = input_171;
      end
      8'b10101100 : begin
        result = input_172;
      end
      8'b10101101 : begin
        result = input_173;
      end
      8'b10101110 : begin
        result = input_174;
      end
      default : begin
        result = input_175;
      end
    endcase
    MUX_v_8_176_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AddRoundKey
// ------------------------------------------------------------------


module AddRoundKey (
  clk, rst_n, round_rsc_dat, round_triosy_lz, state_rsc_zout, state_rsc_lzout, state_rsc_zin,
      state_triosy_lz, RoundKey_rsc_dat, RoundKey_triosy_lz
);
  input clk;
  input rst_n;
  input [7:0] round_rsc_dat;
  output round_triosy_lz;
  output [127:0] state_rsc_zout;
  output state_rsc_lzout;
  input [127:0] state_rsc_zin;
  output state_triosy_lz;
  input [1415:0] RoundKey_rsc_dat;
  output RoundKey_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  AddRoundKey_core AddRoundKey_core_inst (
      .clk(clk),
      .rst_n(rst_n),
      .round_rsc_dat(round_rsc_dat),
      .round_triosy_lz(round_triosy_lz),
      .state_rsc_zout(state_rsc_zout),
      .state_rsc_lzout(state_rsc_lzout),
      .state_rsc_zin(state_rsc_zin),
      .state_triosy_lz(state_triosy_lz),
      .RoundKey_rsc_dat(RoundKey_rsc_dat),
      .RoundKey_triosy_lz(RoundKey_triosy_lz)
    );
endmodule



