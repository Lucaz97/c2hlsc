
//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_inout_prereg_en_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2019 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_inout_prereg_en_v1 (din, ldout, dout, zin, lzout, zout);

    parameter integer rscid = 1;
    parameter integer width = 8;

    output [width-1:0] din;
    input              ldout;
    input  [width-1:0] dout;
    input  [width-1:0] zin;
    output             lzout;
    output [width-1:0] zout;

    wire   [width-1:0] din;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzout = ldout;
    assign din = zin;
    assign zout = dout;

endmodule



//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ../td_ccore_solutions/ROM_1i8_1o8_6cd8ed6ecb89da3c4ea51c9925c1afffbc_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   lc4976@hansolo.poly.edu
//  Generated date: Tue Apr  9 23:32:55 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i8_1o8_6cd8ed6ecb89da3c4ea51c9925c1afffbc
// ------------------------------------------------------------------


module ROM_1i8_1o8_6cd8ed6ecb89da3c4ea51c9925c1afffbc (
  I_1, O_1
);
  input [7:0] I_1;
  output [7:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_8_256_2(8'b01100011, 8'b01111100, 8'b01110111, 8'b01111011,
      8'b11110010, 8'b01101011, 8'b01101111, 8'b11000101, 8'b00110000, 8'b00000001,
      8'b01100111, 8'b00101011, 8'b11111110, 8'b11010111, 8'b10101011, 8'b01110110,
      8'b11001010, 8'b10000010, 8'b11001001, 8'b01111101, 8'b11111010, 8'b01011001,
      8'b01000111, 8'b11110000, 8'b10101101, 8'b11010100, 8'b10100010, 8'b10101111,
      8'b10011100, 8'b10100100, 8'b01110010, 8'b11000000, 8'b10110111, 8'b11111101,
      8'b10010011, 8'b00100110, 8'b00110110, 8'b00111111, 8'b11110111, 8'b11001100,
      8'b00110100, 8'b10100101, 8'b11100101, 8'b11110001, 8'b01110001, 8'b11011000,
      8'b00110001, 8'b00010101, 8'b00000100, 8'b11000111, 8'b00100011, 8'b11000011,
      8'b00011000, 8'b10010110, 8'b00000101, 8'b10011010, 8'b00000111, 8'b00010010,
      8'b10000000, 8'b11100010, 8'b11101011, 8'b00100111, 8'b10110010, 8'b01110101,
      8'b00001001, 8'b10000011, 8'b00101100, 8'b00011010, 8'b00011011, 8'b01101110,
      8'b01011010, 8'b10100000, 8'b01010010, 8'b00111011, 8'b11010110, 8'b10110011,
      8'b00101001, 8'b11100011, 8'b00101111, 8'b10000100, 8'b01010011, 8'b11010001,
      8'b00000000, 8'b11101101, 8'b00100000, 8'b11111100, 8'b10110001, 8'b01011011,
      8'b01101010, 8'b11001011, 8'b10111110, 8'b00111001, 8'b01001010, 8'b01001100,
      8'b01011000, 8'b11001111, 8'b11010000, 8'b11101111, 8'b10101010, 8'b11111011,
      8'b01000011, 8'b01001101, 8'b00110011, 8'b10000101, 8'b01000101, 8'b11111001,
      8'b00000010, 8'b01111111, 8'b01010000, 8'b00111100, 8'b10011111, 8'b10101000,
      8'b01010001, 8'b10100011, 8'b01000000, 8'b10001111, 8'b10010010, 8'b10011101,
      8'b00111000, 8'b11110101, 8'b10111100, 8'b10110110, 8'b11011010, 8'b00100001,
      8'b00010000, 8'b11111111, 8'b11110011, 8'b11010010, 8'b11001101, 8'b00001100,
      8'b00010011, 8'b11101100, 8'b01011111, 8'b10010111, 8'b01000100, 8'b00010111,
      8'b11000100, 8'b10100111, 8'b01111110, 8'b00111101, 8'b01100100, 8'b01011101,
      8'b00011001, 8'b01110011, 8'b01100000, 8'b10000001, 8'b01001111, 8'b11011100,
      8'b00100010, 8'b00101010, 8'b10010000, 8'b10001000, 8'b01000110, 8'b11101110,
      8'b10111000, 8'b00010100, 8'b11011110, 8'b01011110, 8'b00001011, 8'b11011011,
      8'b11100000, 8'b00110010, 8'b00111010, 8'b00001010, 8'b01001001, 8'b00000110,
      8'b00100100, 8'b01011100, 8'b11000010, 8'b11010011, 8'b10101100, 8'b01100010,
      8'b10010001, 8'b10010101, 8'b11100100, 8'b01111001, 8'b11100111, 8'b11001000,
      8'b00110111, 8'b01101101, 8'b10001101, 8'b11010101, 8'b01001110, 8'b10101001,
      8'b01101100, 8'b01010110, 8'b11110100, 8'b11101010, 8'b01100101, 8'b01111010,
      8'b10101110, 8'b00001000, 8'b10111010, 8'b01111000, 8'b00100101, 8'b00101110,
      8'b00011100, 8'b10100110, 8'b10110100, 8'b11000110, 8'b11101000, 8'b11011101,
      8'b01110100, 8'b00011111, 8'b01001011, 8'b10111101, 8'b10001011, 8'b10001010,
      8'b01110000, 8'b00111110, 8'b10110101, 8'b01100110, 8'b01001000, 8'b00000011,
      8'b11110110, 8'b00001110, 8'b01100001, 8'b00110101, 8'b01010111, 8'b10111001,
      8'b10000110, 8'b11000001, 8'b00011101, 8'b10011110, 8'b11100001, 8'b11111000,
      8'b10011000, 8'b00010001, 8'b01101001, 8'b11011001, 8'b10001110, 8'b10010100,
      8'b10011011, 8'b00011110, 8'b10000111, 8'b11101001, 8'b11001110, 8'b01010101,
      8'b00101000, 8'b11011111, 8'b10001100, 8'b10100001, 8'b10001001, 8'b00001101,
      8'b10111111, 8'b11100110, 8'b01000010, 8'b01101000, 8'b01000001, 8'b10011001,
      8'b00101101, 8'b00001111, 8'b10110000, 8'b01010100, 8'b10111011, 8'b00010110,
      I_1);

  function automatic [7:0] MUX_v_8_256_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [7:0] input_16;
    input [7:0] input_17;
    input [7:0] input_18;
    input [7:0] input_19;
    input [7:0] input_20;
    input [7:0] input_21;
    input [7:0] input_22;
    input [7:0] input_23;
    input [7:0] input_24;
    input [7:0] input_25;
    input [7:0] input_26;
    input [7:0] input_27;
    input [7:0] input_28;
    input [7:0] input_29;
    input [7:0] input_30;
    input [7:0] input_31;
    input [7:0] input_32;
    input [7:0] input_33;
    input [7:0] input_34;
    input [7:0] input_35;
    input [7:0] input_36;
    input [7:0] input_37;
    input [7:0] input_38;
    input [7:0] input_39;
    input [7:0] input_40;
    input [7:0] input_41;
    input [7:0] input_42;
    input [7:0] input_43;
    input [7:0] input_44;
    input [7:0] input_45;
    input [7:0] input_46;
    input [7:0] input_47;
    input [7:0] input_48;
    input [7:0] input_49;
    input [7:0] input_50;
    input [7:0] input_51;
    input [7:0] input_52;
    input [7:0] input_53;
    input [7:0] input_54;
    input [7:0] input_55;
    input [7:0] input_56;
    input [7:0] input_57;
    input [7:0] input_58;
    input [7:0] input_59;
    input [7:0] input_60;
    input [7:0] input_61;
    input [7:0] input_62;
    input [7:0] input_63;
    input [7:0] input_64;
    input [7:0] input_65;
    input [7:0] input_66;
    input [7:0] input_67;
    input [7:0] input_68;
    input [7:0] input_69;
    input [7:0] input_70;
    input [7:0] input_71;
    input [7:0] input_72;
    input [7:0] input_73;
    input [7:0] input_74;
    input [7:0] input_75;
    input [7:0] input_76;
    input [7:0] input_77;
    input [7:0] input_78;
    input [7:0] input_79;
    input [7:0] input_80;
    input [7:0] input_81;
    input [7:0] input_82;
    input [7:0] input_83;
    input [7:0] input_84;
    input [7:0] input_85;
    input [7:0] input_86;
    input [7:0] input_87;
    input [7:0] input_88;
    input [7:0] input_89;
    input [7:0] input_90;
    input [7:0] input_91;
    input [7:0] input_92;
    input [7:0] input_93;
    input [7:0] input_94;
    input [7:0] input_95;
    input [7:0] input_96;
    input [7:0] input_97;
    input [7:0] input_98;
    input [7:0] input_99;
    input [7:0] input_100;
    input [7:0] input_101;
    input [7:0] input_102;
    input [7:0] input_103;
    input [7:0] input_104;
    input [7:0] input_105;
    input [7:0] input_106;
    input [7:0] input_107;
    input [7:0] input_108;
    input [7:0] input_109;
    input [7:0] input_110;
    input [7:0] input_111;
    input [7:0] input_112;
    input [7:0] input_113;
    input [7:0] input_114;
    input [7:0] input_115;
    input [7:0] input_116;
    input [7:0] input_117;
    input [7:0] input_118;
    input [7:0] input_119;
    input [7:0] input_120;
    input [7:0] input_121;
    input [7:0] input_122;
    input [7:0] input_123;
    input [7:0] input_124;
    input [7:0] input_125;
    input [7:0] input_126;
    input [7:0] input_127;
    input [7:0] input_128;
    input [7:0] input_129;
    input [7:0] input_130;
    input [7:0] input_131;
    input [7:0] input_132;
    input [7:0] input_133;
    input [7:0] input_134;
    input [7:0] input_135;
    input [7:0] input_136;
    input [7:0] input_137;
    input [7:0] input_138;
    input [7:0] input_139;
    input [7:0] input_140;
    input [7:0] input_141;
    input [7:0] input_142;
    input [7:0] input_143;
    input [7:0] input_144;
    input [7:0] input_145;
    input [7:0] input_146;
    input [7:0] input_147;
    input [7:0] input_148;
    input [7:0] input_149;
    input [7:0] input_150;
    input [7:0] input_151;
    input [7:0] input_152;
    input [7:0] input_153;
    input [7:0] input_154;
    input [7:0] input_155;
    input [7:0] input_156;
    input [7:0] input_157;
    input [7:0] input_158;
    input [7:0] input_159;
    input [7:0] input_160;
    input [7:0] input_161;
    input [7:0] input_162;
    input [7:0] input_163;
    input [7:0] input_164;
    input [7:0] input_165;
    input [7:0] input_166;
    input [7:0] input_167;
    input [7:0] input_168;
    input [7:0] input_169;
    input [7:0] input_170;
    input [7:0] input_171;
    input [7:0] input_172;
    input [7:0] input_173;
    input [7:0] input_174;
    input [7:0] input_175;
    input [7:0] input_176;
    input [7:0] input_177;
    input [7:0] input_178;
    input [7:0] input_179;
    input [7:0] input_180;
    input [7:0] input_181;
    input [7:0] input_182;
    input [7:0] input_183;
    input [7:0] input_184;
    input [7:0] input_185;
    input [7:0] input_186;
    input [7:0] input_187;
    input [7:0] input_188;
    input [7:0] input_189;
    input [7:0] input_190;
    input [7:0] input_191;
    input [7:0] input_192;
    input [7:0] input_193;
    input [7:0] input_194;
    input [7:0] input_195;
    input [7:0] input_196;
    input [7:0] input_197;
    input [7:0] input_198;
    input [7:0] input_199;
    input [7:0] input_200;
    input [7:0] input_201;
    input [7:0] input_202;
    input [7:0] input_203;
    input [7:0] input_204;
    input [7:0] input_205;
    input [7:0] input_206;
    input [7:0] input_207;
    input [7:0] input_208;
    input [7:0] input_209;
    input [7:0] input_210;
    input [7:0] input_211;
    input [7:0] input_212;
    input [7:0] input_213;
    input [7:0] input_214;
    input [7:0] input_215;
    input [7:0] input_216;
    input [7:0] input_217;
    input [7:0] input_218;
    input [7:0] input_219;
    input [7:0] input_220;
    input [7:0] input_221;
    input [7:0] input_222;
    input [7:0] input_223;
    input [7:0] input_224;
    input [7:0] input_225;
    input [7:0] input_226;
    input [7:0] input_227;
    input [7:0] input_228;
    input [7:0] input_229;
    input [7:0] input_230;
    input [7:0] input_231;
    input [7:0] input_232;
    input [7:0] input_233;
    input [7:0] input_234;
    input [7:0] input_235;
    input [7:0] input_236;
    input [7:0] input_237;
    input [7:0] input_238;
    input [7:0] input_239;
    input [7:0] input_240;
    input [7:0] input_241;
    input [7:0] input_242;
    input [7:0] input_243;
    input [7:0] input_244;
    input [7:0] input_245;
    input [7:0] input_246;
    input [7:0] input_247;
    input [7:0] input_248;
    input [7:0] input_249;
    input [7:0] input_250;
    input [7:0] input_251;
    input [7:0] input_252;
    input [7:0] input_253;
    input [7:0] input_254;
    input [7:0] input_255;
    input [7:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      8'b00000000 : begin
        result = input_0;
      end
      8'b00000001 : begin
        result = input_1;
      end
      8'b00000010 : begin
        result = input_2;
      end
      8'b00000011 : begin
        result = input_3;
      end
      8'b00000100 : begin
        result = input_4;
      end
      8'b00000101 : begin
        result = input_5;
      end
      8'b00000110 : begin
        result = input_6;
      end
      8'b00000111 : begin
        result = input_7;
      end
      8'b00001000 : begin
        result = input_8;
      end
      8'b00001001 : begin
        result = input_9;
      end
      8'b00001010 : begin
        result = input_10;
      end
      8'b00001011 : begin
        result = input_11;
      end
      8'b00001100 : begin
        result = input_12;
      end
      8'b00001101 : begin
        result = input_13;
      end
      8'b00001110 : begin
        result = input_14;
      end
      8'b00001111 : begin
        result = input_15;
      end
      8'b00010000 : begin
        result = input_16;
      end
      8'b00010001 : begin
        result = input_17;
      end
      8'b00010010 : begin
        result = input_18;
      end
      8'b00010011 : begin
        result = input_19;
      end
      8'b00010100 : begin
        result = input_20;
      end
      8'b00010101 : begin
        result = input_21;
      end
      8'b00010110 : begin
        result = input_22;
      end
      8'b00010111 : begin
        result = input_23;
      end
      8'b00011000 : begin
        result = input_24;
      end
      8'b00011001 : begin
        result = input_25;
      end
      8'b00011010 : begin
        result = input_26;
      end
      8'b00011011 : begin
        result = input_27;
      end
      8'b00011100 : begin
        result = input_28;
      end
      8'b00011101 : begin
        result = input_29;
      end
      8'b00011110 : begin
        result = input_30;
      end
      8'b00011111 : begin
        result = input_31;
      end
      8'b00100000 : begin
        result = input_32;
      end
      8'b00100001 : begin
        result = input_33;
      end
      8'b00100010 : begin
        result = input_34;
      end
      8'b00100011 : begin
        result = input_35;
      end
      8'b00100100 : begin
        result = input_36;
      end
      8'b00100101 : begin
        result = input_37;
      end
      8'b00100110 : begin
        result = input_38;
      end
      8'b00100111 : begin
        result = input_39;
      end
      8'b00101000 : begin
        result = input_40;
      end
      8'b00101001 : begin
        result = input_41;
      end
      8'b00101010 : begin
        result = input_42;
      end
      8'b00101011 : begin
        result = input_43;
      end
      8'b00101100 : begin
        result = input_44;
      end
      8'b00101101 : begin
        result = input_45;
      end
      8'b00101110 : begin
        result = input_46;
      end
      8'b00101111 : begin
        result = input_47;
      end
      8'b00110000 : begin
        result = input_48;
      end
      8'b00110001 : begin
        result = input_49;
      end
      8'b00110010 : begin
        result = input_50;
      end
      8'b00110011 : begin
        result = input_51;
      end
      8'b00110100 : begin
        result = input_52;
      end
      8'b00110101 : begin
        result = input_53;
      end
      8'b00110110 : begin
        result = input_54;
      end
      8'b00110111 : begin
        result = input_55;
      end
      8'b00111000 : begin
        result = input_56;
      end
      8'b00111001 : begin
        result = input_57;
      end
      8'b00111010 : begin
        result = input_58;
      end
      8'b00111011 : begin
        result = input_59;
      end
      8'b00111100 : begin
        result = input_60;
      end
      8'b00111101 : begin
        result = input_61;
      end
      8'b00111110 : begin
        result = input_62;
      end
      8'b00111111 : begin
        result = input_63;
      end
      8'b01000000 : begin
        result = input_64;
      end
      8'b01000001 : begin
        result = input_65;
      end
      8'b01000010 : begin
        result = input_66;
      end
      8'b01000011 : begin
        result = input_67;
      end
      8'b01000100 : begin
        result = input_68;
      end
      8'b01000101 : begin
        result = input_69;
      end
      8'b01000110 : begin
        result = input_70;
      end
      8'b01000111 : begin
        result = input_71;
      end
      8'b01001000 : begin
        result = input_72;
      end
      8'b01001001 : begin
        result = input_73;
      end
      8'b01001010 : begin
        result = input_74;
      end
      8'b01001011 : begin
        result = input_75;
      end
      8'b01001100 : begin
        result = input_76;
      end
      8'b01001101 : begin
        result = input_77;
      end
      8'b01001110 : begin
        result = input_78;
      end
      8'b01001111 : begin
        result = input_79;
      end
      8'b01010000 : begin
        result = input_80;
      end
      8'b01010001 : begin
        result = input_81;
      end
      8'b01010010 : begin
        result = input_82;
      end
      8'b01010011 : begin
        result = input_83;
      end
      8'b01010100 : begin
        result = input_84;
      end
      8'b01010101 : begin
        result = input_85;
      end
      8'b01010110 : begin
        result = input_86;
      end
      8'b01010111 : begin
        result = input_87;
      end
      8'b01011000 : begin
        result = input_88;
      end
      8'b01011001 : begin
        result = input_89;
      end
      8'b01011010 : begin
        result = input_90;
      end
      8'b01011011 : begin
        result = input_91;
      end
      8'b01011100 : begin
        result = input_92;
      end
      8'b01011101 : begin
        result = input_93;
      end
      8'b01011110 : begin
        result = input_94;
      end
      8'b01011111 : begin
        result = input_95;
      end
      8'b01100000 : begin
        result = input_96;
      end
      8'b01100001 : begin
        result = input_97;
      end
      8'b01100010 : begin
        result = input_98;
      end
      8'b01100011 : begin
        result = input_99;
      end
      8'b01100100 : begin
        result = input_100;
      end
      8'b01100101 : begin
        result = input_101;
      end
      8'b01100110 : begin
        result = input_102;
      end
      8'b01100111 : begin
        result = input_103;
      end
      8'b01101000 : begin
        result = input_104;
      end
      8'b01101001 : begin
        result = input_105;
      end
      8'b01101010 : begin
        result = input_106;
      end
      8'b01101011 : begin
        result = input_107;
      end
      8'b01101100 : begin
        result = input_108;
      end
      8'b01101101 : begin
        result = input_109;
      end
      8'b01101110 : begin
        result = input_110;
      end
      8'b01101111 : begin
        result = input_111;
      end
      8'b01110000 : begin
        result = input_112;
      end
      8'b01110001 : begin
        result = input_113;
      end
      8'b01110010 : begin
        result = input_114;
      end
      8'b01110011 : begin
        result = input_115;
      end
      8'b01110100 : begin
        result = input_116;
      end
      8'b01110101 : begin
        result = input_117;
      end
      8'b01110110 : begin
        result = input_118;
      end
      8'b01110111 : begin
        result = input_119;
      end
      8'b01111000 : begin
        result = input_120;
      end
      8'b01111001 : begin
        result = input_121;
      end
      8'b01111010 : begin
        result = input_122;
      end
      8'b01111011 : begin
        result = input_123;
      end
      8'b01111100 : begin
        result = input_124;
      end
      8'b01111101 : begin
        result = input_125;
      end
      8'b01111110 : begin
        result = input_126;
      end
      8'b01111111 : begin
        result = input_127;
      end
      8'b10000000 : begin
        result = input_128;
      end
      8'b10000001 : begin
        result = input_129;
      end
      8'b10000010 : begin
        result = input_130;
      end
      8'b10000011 : begin
        result = input_131;
      end
      8'b10000100 : begin
        result = input_132;
      end
      8'b10000101 : begin
        result = input_133;
      end
      8'b10000110 : begin
        result = input_134;
      end
      8'b10000111 : begin
        result = input_135;
      end
      8'b10001000 : begin
        result = input_136;
      end
      8'b10001001 : begin
        result = input_137;
      end
      8'b10001010 : begin
        result = input_138;
      end
      8'b10001011 : begin
        result = input_139;
      end
      8'b10001100 : begin
        result = input_140;
      end
      8'b10001101 : begin
        result = input_141;
      end
      8'b10001110 : begin
        result = input_142;
      end
      8'b10001111 : begin
        result = input_143;
      end
      8'b10010000 : begin
        result = input_144;
      end
      8'b10010001 : begin
        result = input_145;
      end
      8'b10010010 : begin
        result = input_146;
      end
      8'b10010011 : begin
        result = input_147;
      end
      8'b10010100 : begin
        result = input_148;
      end
      8'b10010101 : begin
        result = input_149;
      end
      8'b10010110 : begin
        result = input_150;
      end
      8'b10010111 : begin
        result = input_151;
      end
      8'b10011000 : begin
        result = input_152;
      end
      8'b10011001 : begin
        result = input_153;
      end
      8'b10011010 : begin
        result = input_154;
      end
      8'b10011011 : begin
        result = input_155;
      end
      8'b10011100 : begin
        result = input_156;
      end
      8'b10011101 : begin
        result = input_157;
      end
      8'b10011110 : begin
        result = input_158;
      end
      8'b10011111 : begin
        result = input_159;
      end
      8'b10100000 : begin
        result = input_160;
      end
      8'b10100001 : begin
        result = input_161;
      end
      8'b10100010 : begin
        result = input_162;
      end
      8'b10100011 : begin
        result = input_163;
      end
      8'b10100100 : begin
        result = input_164;
      end
      8'b10100101 : begin
        result = input_165;
      end
      8'b10100110 : begin
        result = input_166;
      end
      8'b10100111 : begin
        result = input_167;
      end
      8'b10101000 : begin
        result = input_168;
      end
      8'b10101001 : begin
        result = input_169;
      end
      8'b10101010 : begin
        result = input_170;
      end
      8'b10101011 : begin
        result = input_171;
      end
      8'b10101100 : begin
        result = input_172;
      end
      8'b10101101 : begin
        result = input_173;
      end
      8'b10101110 : begin
        result = input_174;
      end
      8'b10101111 : begin
        result = input_175;
      end
      8'b10110000 : begin
        result = input_176;
      end
      8'b10110001 : begin
        result = input_177;
      end
      8'b10110010 : begin
        result = input_178;
      end
      8'b10110011 : begin
        result = input_179;
      end
      8'b10110100 : begin
        result = input_180;
      end
      8'b10110101 : begin
        result = input_181;
      end
      8'b10110110 : begin
        result = input_182;
      end
      8'b10110111 : begin
        result = input_183;
      end
      8'b10111000 : begin
        result = input_184;
      end
      8'b10111001 : begin
        result = input_185;
      end
      8'b10111010 : begin
        result = input_186;
      end
      8'b10111011 : begin
        result = input_187;
      end
      8'b10111100 : begin
        result = input_188;
      end
      8'b10111101 : begin
        result = input_189;
      end
      8'b10111110 : begin
        result = input_190;
      end
      8'b10111111 : begin
        result = input_191;
      end
      8'b11000000 : begin
        result = input_192;
      end
      8'b11000001 : begin
        result = input_193;
      end
      8'b11000010 : begin
        result = input_194;
      end
      8'b11000011 : begin
        result = input_195;
      end
      8'b11000100 : begin
        result = input_196;
      end
      8'b11000101 : begin
        result = input_197;
      end
      8'b11000110 : begin
        result = input_198;
      end
      8'b11000111 : begin
        result = input_199;
      end
      8'b11001000 : begin
        result = input_200;
      end
      8'b11001001 : begin
        result = input_201;
      end
      8'b11001010 : begin
        result = input_202;
      end
      8'b11001011 : begin
        result = input_203;
      end
      8'b11001100 : begin
        result = input_204;
      end
      8'b11001101 : begin
        result = input_205;
      end
      8'b11001110 : begin
        result = input_206;
      end
      8'b11001111 : begin
        result = input_207;
      end
      8'b11010000 : begin
        result = input_208;
      end
      8'b11010001 : begin
        result = input_209;
      end
      8'b11010010 : begin
        result = input_210;
      end
      8'b11010011 : begin
        result = input_211;
      end
      8'b11010100 : begin
        result = input_212;
      end
      8'b11010101 : begin
        result = input_213;
      end
      8'b11010110 : begin
        result = input_214;
      end
      8'b11010111 : begin
        result = input_215;
      end
      8'b11011000 : begin
        result = input_216;
      end
      8'b11011001 : begin
        result = input_217;
      end
      8'b11011010 : begin
        result = input_218;
      end
      8'b11011011 : begin
        result = input_219;
      end
      8'b11011100 : begin
        result = input_220;
      end
      8'b11011101 : begin
        result = input_221;
      end
      8'b11011110 : begin
        result = input_222;
      end
      8'b11011111 : begin
        result = input_223;
      end
      8'b11100000 : begin
        result = input_224;
      end
      8'b11100001 : begin
        result = input_225;
      end
      8'b11100010 : begin
        result = input_226;
      end
      8'b11100011 : begin
        result = input_227;
      end
      8'b11100100 : begin
        result = input_228;
      end
      8'b11100101 : begin
        result = input_229;
      end
      8'b11100110 : begin
        result = input_230;
      end
      8'b11100111 : begin
        result = input_231;
      end
      8'b11101000 : begin
        result = input_232;
      end
      8'b11101001 : begin
        result = input_233;
      end
      8'b11101010 : begin
        result = input_234;
      end
      8'b11101011 : begin
        result = input_235;
      end
      8'b11101100 : begin
        result = input_236;
      end
      8'b11101101 : begin
        result = input_237;
      end
      8'b11101110 : begin
        result = input_238;
      end
      8'b11101111 : begin
        result = input_239;
      end
      8'b11110000 : begin
        result = input_240;
      end
      8'b11110001 : begin
        result = input_241;
      end
      8'b11110010 : begin
        result = input_242;
      end
      8'b11110011 : begin
        result = input_243;
      end
      8'b11110100 : begin
        result = input_244;
      end
      8'b11110101 : begin
        result = input_245;
      end
      8'b11110110 : begin
        result = input_246;
      end
      8'b11110111 : begin
        result = input_247;
      end
      8'b11111000 : begin
        result = input_248;
      end
      8'b11111001 : begin
        result = input_249;
      end
      8'b11111010 : begin
        result = input_250;
      end
      8'b11111011 : begin
        result = input_251;
      end
      8'b11111100 : begin
        result = input_252;
      end
      8'b11111101 : begin
        result = input_253;
      end
      8'b11111110 : begin
        result = input_254;
      end
      default : begin
        result = input_255;
      end
    endcase
    MUX_v_8_256_2 = result;
  end
  endfunction

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   lc4976@hansolo.poly.edu
//  Generated date: Tue Apr  9 23:33:06 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SubBytes_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module SubBytes_core_core_fsm (
  clk, rst_n, fsm_output, for_for_C_1_tr0, for_C_0_tr0
);
  input clk;
  input rst_n;
  output [4:0] fsm_output;
  reg [4:0] fsm_output;
  input for_for_C_1_tr0;
  input for_C_0_tr0;


  // FSM State Type Declaration for SubBytes_core_core_fsm_1
  parameter
    main_C_0 = 3'd0,
    for_for_C_0 = 3'd1,
    for_for_C_1 = 3'd2,
    for_C_0 = 3'd3,
    main_C_1 = 3'd4;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SubBytes_core_core_fsm_1
    case (state_var)
      for_for_C_0 : begin
        fsm_output = 5'b00010;
        state_var_NS = for_for_C_1;
      end
      for_for_C_1 : begin
        fsm_output = 5'b00100;
        if ( for_for_C_1_tr0 ) begin
          state_var_NS = for_C_0;
        end
        else begin
          state_var_NS = for_for_C_0;
        end
      end
      for_C_0 : begin
        fsm_output = 5'b01000;
        if ( for_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 5'b10000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 5'b00001;
        state_var_NS = for_for_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SubBytes_core
// ------------------------------------------------------------------


module SubBytes_core (
  clk, rst_n, state_rsc_zout, state_rsc_lzout, state_rsc_zin, state_triosy_lz
);
  input clk;
  input rst_n;
  output [127:0] state_rsc_zout;
  output state_rsc_lzout;
  input [127:0] state_rsc_zin;
  output state_triosy_lz;


  // Interconnect Declarations
  wire [127:0] state_rsci_din;
  reg state_triosy_obj_ld;
  wire [4:0] fsm_output;
  wire or_dcpl_2;
  wire or_dcpl_3;
  wire or_dcpl_5;
  wire or_dcpl_7;
  wire or_dcpl_9;
  wire or_dcpl_10;
  wire or_dcpl_15;
  wire or_dcpl_20;
  reg [1:0] i_2_0_sva_1_0;
  reg [1:0] j_2_0_sva_1_0;
  wire i_or_cse;
  wire [2:0] z_out;
  wire [3:0] nl_z_out;
  wire [7:0] ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1;

  wire i_not_1_nl;
  wire i_not_nl;
  wire[1:0] for_for_mux_18_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_state_rsci_ldout;
  assign nl_state_rsci_ldout = fsm_output[1];
  wire[7:0] for_for_mux_15_nl;
  wire or_25_nl;
  wire[7:0] for_for_mux_14_nl;
  wire or_24_nl;
  wire[7:0] for_for_mux_13_nl;
  wire or_23_nl;
  wire[7:0] for_for_mux_12_nl;
  wire or_22_nl;
  wire[7:0] for_for_mux_11_nl;
  wire or_20_nl;
  wire[7:0] for_for_mux_10_nl;
  wire or_19_nl;
  wire[7:0] for_for_mux_9_nl;
  wire or_18_nl;
  wire[7:0] for_for_mux_8_nl;
  wire or_17_nl;
  wire[7:0] for_for_mux_7_nl;
  wire or_15_nl;
  wire[7:0] for_for_mux_6_nl;
  wire or_14_nl;
  wire[7:0] for_for_mux_5_nl;
  wire or_13_nl;
  wire[7:0] for_for_mux_4_nl;
  wire or_12_nl;
  wire[7:0] for_for_mux_3_nl;
  wire or_9_nl;
  wire[7:0] for_for_mux_2_nl;
  wire or_7_nl;
  wire[7:0] for_for_mux_1_nl;
  wire or_5_nl;
  wire[7:0] for_for_mux_nl;
  wire for_for_nor_nl;
  wire [127:0] nl_state_rsci_dout;
  assign or_25_nl = or_dcpl_20 | or_dcpl_7;
  assign for_for_mux_15_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[127:120]), or_25_nl);
  assign or_24_nl = or_dcpl_20 | or_dcpl_5;
  assign for_for_mux_14_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[119:112]), or_24_nl);
  assign or_23_nl = or_dcpl_20 | or_dcpl_2;
  assign for_for_mux_13_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[111:104]), or_23_nl);
  assign or_22_nl = or_dcpl_20 | or_dcpl_9;
  assign for_for_mux_12_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[103:96]), or_22_nl);
  assign or_20_nl = or_dcpl_15 | or_dcpl_7;
  assign for_for_mux_11_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[95:88]), or_20_nl);
  assign or_19_nl = or_dcpl_15 | or_dcpl_5;
  assign for_for_mux_10_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[87:80]), or_19_nl);
  assign or_18_nl = or_dcpl_15 | or_dcpl_2;
  assign for_for_mux_9_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[79:72]), or_18_nl);
  assign or_17_nl = or_dcpl_15 | or_dcpl_9;
  assign for_for_mux_8_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[71:64]), or_17_nl);
  assign or_15_nl = or_dcpl_10 | or_dcpl_7;
  assign for_for_mux_7_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[63:56]), or_15_nl);
  assign or_14_nl = or_dcpl_10 | or_dcpl_5;
  assign for_for_mux_6_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[55:48]), or_14_nl);
  assign or_13_nl = or_dcpl_10 | or_dcpl_2;
  assign for_for_mux_5_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[47:40]), or_13_nl);
  assign or_12_nl = or_dcpl_10 | or_dcpl_9;
  assign for_for_mux_4_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[39:32]), or_12_nl);
  assign or_9_nl = or_dcpl_3 | or_dcpl_7;
  assign for_for_mux_3_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[31:24]), or_9_nl);
  assign or_7_nl = or_dcpl_3 | or_dcpl_5;
  assign for_for_mux_2_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[23:16]), or_7_nl);
  assign or_5_nl = or_dcpl_3 | or_dcpl_2;
  assign for_for_mux_1_nl = MUX_v_8_2_2(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      (state_rsci_din[15:8]), or_5_nl);
  assign for_for_nor_nl = ~(((i_2_0_sva_1_0[0]) & (~((j_2_0_sva_1_0!=2'b00) | (i_2_0_sva_1_0[1]))))
      | ((i_2_0_sva_1_0[1]) & (~((j_2_0_sva_1_0!=2'b00) | (i_2_0_sva_1_0[0])))) |
      ((i_2_0_sva_1_0==2'b11) & (j_2_0_sva_1_0==2'b00)) | ((j_2_0_sva_1_0[0]) & (~((j_2_0_sva_1_0[1])
      | (i_2_0_sva_1_0!=2'b00)))) | ((j_2_0_sva_1_0[0]) & (i_2_0_sva_1_0[0]) & (~((j_2_0_sva_1_0[1])
      | (i_2_0_sva_1_0[1])))) | ((j_2_0_sva_1_0[0]) & (i_2_0_sva_1_0[1]) & (~((j_2_0_sva_1_0[1])
      | (i_2_0_sva_1_0[0])))) | ((j_2_0_sva_1_0[0]) & (i_2_0_sva_1_0==2'b11) & (~
      (j_2_0_sva_1_0[1]))) | ((j_2_0_sva_1_0[1]) & (~((j_2_0_sva_1_0[0]) | (i_2_0_sva_1_0!=2'b00))))
      | ((j_2_0_sva_1_0[1]) & (i_2_0_sva_1_0[0]) & (~((j_2_0_sva_1_0[0]) | (i_2_0_sva_1_0[1]))))
      | ((j_2_0_sva_1_0[1]) & (i_2_0_sva_1_0[1]) & (~((j_2_0_sva_1_0[0]) | (i_2_0_sva_1_0[0]))))
      | ((j_2_0_sva_1_0[1]) & (i_2_0_sva_1_0==2'b11) & (~ (j_2_0_sva_1_0[0]))) |
      ((j_2_0_sva_1_0==2'b11) & (i_2_0_sva_1_0==2'b00)) | ((j_2_0_sva_1_0==2'b11)
      & (i_2_0_sva_1_0==2'b01)) | ((j_2_0_sva_1_0==2'b11) & (i_2_0_sva_1_0==2'b10))
      | ((j_2_0_sva_1_0==2'b11) & (i_2_0_sva_1_0==2'b11)));
  assign for_for_mux_nl = MUX_v_8_2_2((state_rsci_din[7:0]), ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1,
      for_for_nor_nl);
  assign nl_state_rsci_dout = {for_for_mux_15_nl , for_for_mux_14_nl , for_for_mux_13_nl
      , for_for_mux_12_nl , for_for_mux_11_nl , for_for_mux_10_nl , for_for_mux_9_nl
      , for_for_mux_8_nl , for_for_mux_7_nl , for_for_mux_6_nl , for_for_mux_5_nl
      , for_for_mux_4_nl , for_for_mux_3_nl , for_for_mux_2_nl , for_for_mux_1_nl
      , for_for_mux_nl};
  wire [7:0] nl_U_ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_rg_I_1;
  assign nl_U_ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_rg_I_1 = MUX_v_8_16_2((state_rsci_din[7:0]),
      (state_rsci_din[15:8]), (state_rsci_din[23:16]), (state_rsci_din[31:24]), (state_rsci_din[39:32]),
      (state_rsci_din[47:40]), (state_rsci_din[55:48]), (state_rsci_din[63:56]),
      (state_rsci_din[71:64]), (state_rsci_din[79:72]), (state_rsci_din[87:80]),
      (state_rsci_din[95:88]), (state_rsci_din[103:96]), (state_rsci_din[111:104]),
      (state_rsci_din[119:112]), (state_rsci_din[127:120]), {j_2_0_sva_1_0 , i_2_0_sva_1_0});
  wire  nl_SubBytes_core_core_fsm_inst_for_for_C_1_tr0;
  assign nl_SubBytes_core_core_fsm_inst_for_for_C_1_tr0 = z_out[2];
  wire  nl_SubBytes_core_core_fsm_inst_for_C_0_tr0;
  assign nl_SubBytes_core_core_fsm_inst_for_C_0_tr0 = z_out[2];
  mgc_inout_prereg_en_v1 #(.rscid(32'sd1),
  .width(32'sd128)) state_rsci (
      .din(state_rsci_din),
      .ldout(nl_state_rsci_ldout),
      .dout(nl_state_rsci_dout[127:0]),
      .zin(state_rsc_zin),
      .lzout(state_rsc_lzout),
      .zout(state_rsc_zout)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) state_triosy_obj (
      .ld(state_triosy_obj_ld),
      .lz(state_triosy_lz)
    );
  ROM_1i8_1o8_6cd8ed6ecb89da3c4ea51c9925c1afffbc  U_ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_rg
      (
      .I_1(nl_U_ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_rg_I_1[7:0]),
      .O_1(ROM_1i8_1o8_ec965ae3708891513d2041cf4eab49d42f_1)
    );
  SubBytes_core_core_fsm SubBytes_core_core_fsm_inst (
      .clk(clk),
      .rst_n(rst_n),
      .fsm_output(fsm_output),
      .for_for_C_1_tr0(nl_SubBytes_core_core_fsm_inst_for_for_C_1_tr0),
      .for_C_0_tr0(nl_SubBytes_core_core_fsm_inst_for_C_0_tr0)
    );
  assign i_or_cse = (fsm_output[0]) | (fsm_output[3]);
  assign or_dcpl_2 = (i_2_0_sva_1_0!=2'b01);
  assign or_dcpl_3 = (j_2_0_sva_1_0!=2'b00);
  assign or_dcpl_5 = (i_2_0_sva_1_0!=2'b10);
  assign or_dcpl_7 = ~((i_2_0_sva_1_0==2'b11));
  assign or_dcpl_9 = (i_2_0_sva_1_0!=2'b00);
  assign or_dcpl_10 = (j_2_0_sva_1_0!=2'b01);
  assign or_dcpl_15 = (j_2_0_sva_1_0!=2'b10);
  assign or_dcpl_20 = ~((j_2_0_sva_1_0==2'b11));
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      i_2_0_sva_1_0 <= 2'b00;
    end
    else if ( i_or_cse ) begin
      i_2_0_sva_1_0 <= MUX_v_2_2_2(2'b00, (z_out[1:0]), i_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      j_2_0_sva_1_0 <= 2'b00;
    end
    else if ( (fsm_output[2]) | i_or_cse ) begin
      j_2_0_sva_1_0 <= MUX_v_2_2_2(2'b00, (z_out[1:0]), i_not_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      state_triosy_obj_ld <= 1'b0;
    end
    else begin
      state_triosy_obj_ld <= (z_out[2]) & (fsm_output[3]);
    end
  end
  assign i_not_1_nl = ~ (fsm_output[0]);
  assign i_not_nl = ~ i_or_cse;
  assign for_for_mux_18_nl = MUX_v_2_2_2(j_2_0_sva_1_0, i_2_0_sva_1_0, fsm_output[3]);
  assign nl_z_out = conv_u2u_2_3(for_for_mux_18_nl) + 3'b001;
  assign z_out = nl_z_out[2:0];

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_16_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [3:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_8_16_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SubBytes
// ------------------------------------------------------------------


module SubBytes (
  clk, rst_n, state_rsc_zout, state_rsc_lzout, state_rsc_zin, state_triosy_lz
);
  input clk;
  input rst_n;
  output [127:0] state_rsc_zout;
  output state_rsc_lzout;
  input [127:0] state_rsc_zin;
  output state_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  SubBytes_core SubBytes_core_inst (
      .clk(clk),
      .rst_n(rst_n),
      .state_rsc_zout(state_rsc_zout),
      .state_rsc_lzout(state_rsc_lzout),
      .state_rsc_zin(state_rsc_zin),
      .state_triosy_lz(state_triosy_lz)
    );
endmodule



